// Benchmark "sin" written by ABC on Fri Feb  7 13:41:11 2014

module sin ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63;
  wire n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
    n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843;
  bufx g0000(.A(n2818), .O(po00));
  bufx g0001(.A(n2817), .O(po01));
  bufx g0002(.A(n2816), .O(po02));
  bufx g0003(.A(n2815), .O(po03));
  bufx g0004(.A(n2814), .O(po04));
  bufx g0005(.A(n2813), .O(po05));
  bufx g0006(.A(n2812), .O(po06));
  bufx g0007(.A(n2811), .O(po07));
  bufx g0008(.A(n2810), .O(po08));
  bufx g0009(.A(n2809), .O(po09));
  bufx g0010(.A(n2808), .O(po10));
  bufx g0011(.A(n2807), .O(po11));
  bufx g0012(.A(n2806), .O(po12));
  bufx g0013(.A(n2805), .O(po13));
  bufx g0014(.A(n2804), .O(po14));
  bufx g0015(.A(n2803), .O(po15));
  bufx g0016(.A(n2802), .O(po16));
  bufx g0017(.A(n2801), .O(po17));
  bufx g0018(.A(n2800), .O(po18));
  bufx g0019(.A(n2799), .O(po19));
  bufx g0020(.A(n2798), .O(po20));
  bufx g0021(.A(n2797), .O(po21));
  bufx g0022(.A(n2796), .O(po22));
  bufx g0023(.A(n2795), .O(po23));
  bufx g0024(.A(n2794), .O(po24));
  bufx g0025(.A(n2793), .O(po25));
  bufx g0026(.A(n2792), .O(po26));
  bufx g0027(.A(n2791), .O(po27));
  bufx g0028(.A(n2790), .O(po28));
  bufx g0029(.A(n2789), .O(po29));
  bufx g0030(.A(n2788), .O(po30));
  bufx g0031(.A(n2787), .O(po31));
  bufx g0032(.A(n2786), .O(po32));
  bufx g0033(.A(n2785), .O(po33));
  bufx g0034(.A(n2784), .O(po34));
  bufx g0035(.A(n2783), .O(po35));
  bufx g0036(.A(n2782), .O(po36));
  bufx g0037(.A(n2781), .O(po37));
  bufx g0038(.A(n2780), .O(po38));
  bufx g0039(.A(n2779), .O(po39));
  bufx g0040(.A(n2778), .O(po40));
  bufx g0041(.A(n2777), .O(po41));
  bufx g0042(.A(n2776), .O(po42));
  bufx g0043(.A(n2775), .O(po43));
  bufx g0044(.A(n2774), .O(po44));
  bufx g0045(.A(n2773), .O(po45));
  bufx g0046(.A(n2772), .O(po46));
  bufx g0047(.A(n2771), .O(po47));
  bufx g0048(.A(n2770), .O(po48));
  bufx g0049(.A(n2769), .O(po49));
  bufx g0050(.A(n2768), .O(po50));
  bufx g0051(.A(n2767), .O(po51));
  bufx g0052(.A(n2742), .O(po52));
  bufx g0053(.A(n2741), .O(po53));
  bufx g0054(.A(n2740), .O(po54));
  bufx g0055(.A(n2739), .O(po55));
  bufx g0056(.A(n2739), .O(po56));
  bufx g0057(.A(n2739), .O(po57));
  bufx g0058(.A(n2739), .O(po58));
  bufx g0059(.A(n2739), .O(po59));
  bufx g0060(.A(n2739), .O(po60));
  bufx g0061(.A(n2739), .O(po61));
  bufx g0062(.A(n2739), .O(po62));
  bufx g0063(.A(n2732), .O(po63));
  orx  g0064(.A(pi03), .B(pi01), .O(n163));
  orx  g0065(.A(pi02), .B(n2354), .O(n164));
  orx  g0066(.A(n2377), .B(n2672), .O(n165));
  andx g0067(.A(n217), .B(n2563), .O(n166));
  orx  g0068(.A(n183), .B(n2485), .O(n167));
  andx g0069(.A(n167), .B(pi05), .O(n168));
  orx  g0070(.A(n2702), .B(n2442), .O(n169));
  andx g0071(.A(n2639), .B(pi00), .O(n170));
  andx g0072(.A(n2602), .B(n2542), .O(n171));
  orx  g0073(.A(n2387), .B(pi03), .O(n172));
  andx g0074(.A(n172), .B(pi05), .O(n173));
  andx g0075(.A(n2675), .B(n2351), .O(n174));
  orx  g0076(.A(n2664), .B(n2378), .O(n175));
  orx  g0077(.A(n2672), .B(n2338), .O(n176));
  andx g0078(.A(n2628), .B(pi00), .O(n177));
  andx g0079(.A(n2650), .B(pi00), .O(n178));
  andx g0080(.A(n2606), .B(n2542), .O(n179));
  andx g0081(.A(pi04), .B(n198), .O(n180));
  orx  g0082(.A(n2355), .B(n2358), .O(n181));
  orx  g0083(.A(n2373), .B(n2757), .O(n182));
  orx  g0084(.A(pi01), .B(pi02), .O(n183));
  orx  g0085(.A(n2463), .B(n2385), .O(n184));
  orx  g0086(.A(pi03), .B(n2357), .O(n185));
  orx  g0087(.A(pi03), .B(n2339), .O(n186));
  orx  g0088(.A(n2384), .B(n2660), .O(n187));
  orx  g0089(.A(pi05), .B(n2660), .O(n188));
  orx  g0090(.A(n2454), .B(n2727), .O(n189));
  orx  g0091(.A(n2338), .B(n2668), .O(n190));
  orx  g0092(.A(pi03), .B(n2397), .O(n191));
  orx  g0093(.A(n2699), .B(n2668), .O(n192));
  orx  g0094(.A(n2398), .B(n2660), .O(n193));
  orx  g0095(.A(n2727), .B(n2660), .O(n194));
  orx  g0096(.A(pi05), .B(n194), .O(n195));
  orx  g0097(.A(pi03), .B(n2372), .O(n196));
  orx  g0098(.A(pi03), .B(n2369), .O(n197));
  orx  g0099(.A(pi03), .B(n2370), .O(n198));
  orx  g0100(.A(pi01), .B(n2486), .O(n199));
  orx  g0101(.A(pi03), .B(n2393), .O(n200));
  orx  g0102(.A(n2664), .B(n2391), .O(n201));
  orx  g0103(.A(pi03), .B(n2330), .O(n202));
  orx  g0104(.A(n2339), .B(n2486), .O(n203));
  orx  g0105(.A(pi05), .B(n2636), .O(n204));
  orx  g0106(.A(n2609), .B(n2370), .O(n205));
  orx  g0107(.A(pi03), .B(n2377), .O(n206));
  orx  g0108(.A(n376), .B(n377), .O(n207));
  orx  g0109(.A(n364), .B(n365), .O(n208));
  orx  g0110(.A(n450), .B(n451), .O(n209));
  orx  g0111(.A(n474), .B(n475), .O(n210));
  orx  g0112(.A(n829), .B(n830), .O(n211));
  orx  g0113(.A(n351), .B(n352), .O(n212));
  andx g0114(.A(n353), .B(n2542), .O(n213));
  orx  g0115(.A(n335), .B(n336), .O(n214));
  orx  g0116(.A(n341), .B(n342), .O(n215));
  orx  g0117(.A(n361), .B(n360), .O(n216));
  orx  g0118(.A(n386), .B(n387), .O(n217));
  orx  g0119(.A(n390), .B(n391), .O(n218));
  orx  g0120(.A(n378), .B(n379), .O(n219));
  andx g0121(.A(pi02), .B(pi03), .O(n220));
  orx  g0122(.A(n366), .B(n367), .O(n221));
  andx g0123(.A(n393), .B(n389), .O(n222));
  orx  g0124(.A(n395), .B(n394), .O(n223));
  orx  g0125(.A(n418), .B(n419), .O(n224));
  orx  g0126(.A(n410), .B(n411), .O(n225));
  orx  g0127(.A(n404), .B(n405), .O(n226));
  orx  g0128(.A(n402), .B(n403), .O(n227));
  orx  g0129(.A(n398), .B(n399), .O(n228));
  orx  g0130(.A(n396), .B(n397), .O(n229));
  andx g0131(.A(n331), .B(n421), .O(n230));
  orx  g0132(.A(n423), .B(n422), .O(n231));
  andx g0133(.A(n452), .B(n2543), .O(n232));
  orx  g0134(.A(n440), .B(n441), .O(n233));
  orx  g0135(.A(n432), .B(n433), .O(n234));
  orx  g0136(.A(n430), .B(n431), .O(n235));
  orx  g0137(.A(n426), .B(n427), .O(n236));
  orx  g0138(.A(n424), .B(n425), .O(n237));
  orx  g0139(.A(n456), .B(n455), .O(n238));
  orx  g0140(.A(n465), .B(n466), .O(n239));
  orx  g0141(.A(n2369), .B(n2672), .O(n240));
  orx  g0142(.A(n2378), .B(n2486), .O(n241));
  andx g0143(.A(n477), .B(n473), .O(n242));
  orx  g0144(.A(n479), .B(n478), .O(n243));
  orx  g0145(.A(n499), .B(n500), .O(n244));
  andx g0146(.A(n2369), .B(n203), .O(n245));
  andx g0147(.A(n502), .B(n2542), .O(n246));
  orx  g0148(.A(n504), .B(n503), .O(n247));
  orx  g0149(.A(n525), .B(n526), .O(n248));
  orx  g0150(.A(n515), .B(n516), .O(n249));
  andx g0151(.A(n529), .B(n2543), .O(n250));
  orx  g0152(.A(n531), .B(n530), .O(n251));
  andx g0153(.A(n2664), .B(n2335), .O(n252));
  andx g0154(.A(n539), .B(n538), .O(n253));
  andx g0155(.A(n2644), .B(n2336), .O(n254));
  andx g0156(.A(n532), .B(n1087), .O(n255));
  orx  g0157(.A(n547), .B(n548), .O(n256));
  orx  g0158(.A(n569), .B(n570), .O(n257));
  andx g0159(.A(n571), .B(n2543), .O(n258));
  orx  g0160(.A(n573), .B(n572), .O(n259));
  andx g0161(.A(n595), .B(n2554), .O(n260));
  orx  g0162(.A(n587), .B(n588), .O(n261));
  orx  g0163(.A(n582), .B(n583), .O(n262));
  orx  g0164(.A(n602), .B(n601), .O(n263));
  andx g0165(.A(n622), .B(n2543), .O(n264));
  orx  g0166(.A(n624), .B(n623), .O(n265));
  orx  g0167(.A(n647), .B(n648), .O(n266));
  orx  g0168(.A(n643), .B(n644), .O(n267));
  andx g0169(.A(n646), .B(n2544), .O(n268));
  orx  g0170(.A(n635), .B(n636), .O(n269));
  orx  g0171(.A(n656), .B(n655), .O(n270));
  andx g0172(.A(n675), .B(n2544), .O(n271));
  orx  g0173(.A(n661), .B(n662), .O(n272));
  orx  g0174(.A(n682), .B(n681), .O(n273));
  orx  g0175(.A(n702), .B(n703), .O(n274));
  andx g0176(.A(n704), .B(n2544), .O(n275));
  orx  g0177(.A(n688), .B(n689), .O(n276));
  orx  g0178(.A(n686), .B(n687), .O(n277));
  orx  g0179(.A(n710), .B(n709), .O(n278));
  orx  g0180(.A(n730), .B(n731), .O(n279));
  orx  g0181(.A(n728), .B(n729), .O(n280));
  andx g0182(.A(n732), .B(n2545), .O(n281));
  orx  g0183(.A(n738), .B(n737), .O(n282));
  orx  g0184(.A(n749), .B(n750), .O(n283));
  orx  g0185(.A(n745), .B(n746), .O(n284));
  andx g0186(.A(n757), .B(n2544), .O(n285));
  orx  g0187(.A(n759), .B(n758), .O(n286));
  andx g0188(.A(n332), .B(n189), .O(n287));
  orx  g0189(.A(n766), .B(n767), .O(n288));
  orx  g0190(.A(n782), .B(n781), .O(n289));
  andx g0191(.A(n798), .B(n2545), .O(n290));
  andx g0192(.A(pi03), .B(n2370), .O(n291));
  orx  g0193(.A(n804), .B(n803), .O(n292));
  andx g0194(.A(n822), .B(n2546), .O(n293));
  orx  g0195(.A(n805), .B(n806), .O(n294));
  orx  g0196(.A(n828), .B(n827), .O(n295));
  andx g0197(.A(n1090), .B(n163), .O(n296));
  andx g0198(.A(n845), .B(n2545), .O(n297));
  orx  g0199(.A(n847), .B(n846), .O(n298));
  orx  g0200(.A(n863), .B(n864), .O(n299));
  andx g0201(.A(n867), .B(n2545), .O(n300));
  orx  g0202(.A(n869), .B(n868), .O(n301));
  andx g0203(.A(n1092), .B(n1081), .O(n302));
  andx g0204(.A(n883), .B(n2546), .O(n303));
  orx  g0205(.A(n885), .B(n884), .O(n304));
  andx g0206(.A(n896), .B(n2546), .O(n305));
  andx g0207(.A(n1093), .B(n194), .O(n306));
  orx  g0208(.A(n902), .B(n901), .O(n307));
  orx  g0209(.A(n922), .B(n921), .O(n308));
  andx g0210(.A(n937), .B(n2546), .O(n309));
  andx g0211(.A(n2597), .B(n1094), .O(n310));
  orx  g0212(.A(n941), .B(n940), .O(n311));
  andx g0213(.A(n960), .B(n958), .O(n312));
  orx  g0214(.A(n962), .B(n961), .O(n313));
  andx g0215(.A(n981), .B(n2547), .O(n314));
  orx  g0216(.A(n963), .B(n964), .O(n315));
  orx  g0217(.A(n985), .B(n984), .O(n316));
  andx g0218(.A(n1001), .B(n2547), .O(n317));
  orx  g0219(.A(n1003), .B(n1002), .O(n318));
  andx g0220(.A(n1020), .B(n2547), .O(n319));
  orx  g0221(.A(n1022), .B(n1021), .O(n320));
  andx g0222(.A(n1041), .B(n2548), .O(n321));
  orx  g0223(.A(n1043), .B(n1042), .O(n322));
  andx g0224(.A(n1058), .B(n2547), .O(n323));
  orx  g0225(.A(n1060), .B(n1059), .O(n324));
  andx g0226(.A(n1077), .B(n2548), .O(n325));
  orx  g0227(.A(n1079), .B(n1078), .O(n326));
  orx  g0228(.A(pi03), .B(n2348), .O(n327));
  orx  g0229(.A(pi02), .B(pi03), .O(n328));
  orx  g0230(.A(pi05), .B(n167), .O(n329));
  orx  g0231(.A(pi05), .B(n198), .O(n330));
  andx g0232(.A(n1080), .B(n2549), .O(n331));
  andx g0233(.A(n2397), .B(n2548), .O(n332));
  andx g0234(.A(n163), .B(n2548), .O(n333));
  andx g0235(.A(n2730), .B(pi05), .O(n334));
  andx g0236(.A(pi03), .B(n2764), .O(n335));
  andx g0237(.A(pi01), .B(n2459), .O(n336));
  andx g0238(.A(n214), .B(n2549), .O(n337));
  andx g0239(.A(n2675), .B(pi05), .O(n338));
  andx g0240(.A(n1098), .B(n2411), .O(n339));
  andx g0241(.A(n1099), .B(pi00), .O(n340));
  andx g0242(.A(n2348), .B(n2460), .O(n341));
  andx g0243(.A(n2394), .B(pi03), .O(n342));
  andx g0244(.A(n1082), .B(n2549), .O(n343));
  andx g0245(.A(n215), .B(pi05), .O(n344));
  andx g0246(.A(n214), .B(pi05), .O(n345));
  andx g0247(.A(n165), .B(n2549), .O(n346));
  andx g0248(.A(n1101), .B(n2427), .O(n347));
  andx g0249(.A(n1102), .B(pi00), .O(n348));
  andx g0250(.A(n1100), .B(n2516), .O(n349));
  andx g0251(.A(n1103), .B(pi04), .O(n350));
  andx g0252(.A(pi03), .B(n2760), .O(n351));
  andx g0253(.A(n2386), .B(n2459), .O(n352));
  andx g0254(.A(n1106), .B(n1105), .O(n353));
  orx  g0255(.A(pi05), .B(n2386), .O(n354));
  orx  g0256(.A(pi05), .B(n185), .O(n355));
  andx g0257(.A(n2731), .B(n2427), .O(n356));
  andx g0258(.A(n2722), .B(pi00), .O(n357));
  andx g0259(.A(n213), .B(n2503), .O(n358));
  andx g0260(.A(n1107), .B(pi04), .O(n359));
  andx g0261(.A(n1104), .B(n2350), .O(n360));
  andx g0262(.A(n1108), .B(pi06), .O(n361));
  andx g0263(.A(n2604), .B(n2550), .O(n362));
  andx g0264(.A(n2603), .B(pi05), .O(n363));
  andx g0265(.A(n2373), .B(pi03), .O(n364));
  andx g0266(.A(n2385), .B(n2474), .O(n365));
  andx g0267(.A(pi01), .B(pi03), .O(n366));
  andx g0268(.A(pi02), .B(n2460), .O(n367));
  andx g0269(.A(n2656), .B(n2550), .O(n368));
  andx g0270(.A(n221), .B(pi05), .O(n369));
  andx g0271(.A(n1109), .B(n2427), .O(n370));
  andx g0272(.A(n1110), .B(pi00), .O(n371));
  andx g0273(.A(n2339), .B(pi03), .O(n372));
  andx g0274(.A(n2384), .B(n2466), .O(n373));
  andx g0275(.A(n1112), .B(n2550), .O(n374));
  andx g0276(.A(n220), .B(pi05), .O(n375));
  andx g0277(.A(pi01), .B(n2361), .O(n376));
  andx g0278(.A(pi02), .B(n2355), .O(n377));
  andx g0279(.A(pi03), .B(n2354), .O(n378));
  andx g0280(.A(n2395), .B(n2460), .O(n379));
  andx g0281(.A(n2368), .B(n2551), .O(n380));
  andx g0282(.A(n219), .B(pi05), .O(n381));
  andx g0283(.A(n1113), .B(n2427), .O(n382));
  andx g0284(.A(n1114), .B(pi00), .O(n383));
  andx g0285(.A(n1111), .B(n2504), .O(n384));
  andx g0286(.A(n1115), .B(pi04), .O(n385));
  andx g0287(.A(n2378), .B(pi03), .O(n386));
  andx g0288(.A(n207), .B(n2461), .O(n387));
  orx  g0289(.A(n166), .B(n2443), .O(n388));
  andx g0290(.A(n1118), .B(n1117), .O(n389));
  andx g0291(.A(n2372), .B(pi03), .O(n390));
  andx g0292(.A(n2393), .B(n2475), .O(n391));
  andx g0293(.A(n1120), .B(n1119), .O(n392));
  andx g0294(.A(n1122), .B(n1121), .O(n393));
  andx g0295(.A(n1116), .B(n2353), .O(n394));
  andx g0296(.A(n222), .B(pi06), .O(n395));
  andx g0297(.A(pi02), .B(pi03), .O(n396));
  andx g0298(.A(n2383), .B(n2461), .O(n397));
  andx g0299(.A(n2370), .B(n2462), .O(n398));
  andx g0300(.A(n2378), .B(pi03), .O(n399));
  andx g0301(.A(n229), .B(n2550), .O(n400));
  andx g0302(.A(n228), .B(pi05), .O(n401));
  andx g0303(.A(n2484), .B(n2359), .O(n402));
  andx g0304(.A(pi03), .B(n2347), .O(n403));
  andx g0305(.A(pi03), .B(n2354), .O(n404));
  andx g0306(.A(n2373), .B(n2462), .O(n405));
  andx g0307(.A(n227), .B(n2551), .O(n406));
  andx g0308(.A(n226), .B(pi05), .O(n407));
  andx g0309(.A(n1123), .B(n2426), .O(n408));
  andx g0310(.A(n1124), .B(pi00), .O(n409));
  andx g0311(.A(n2338), .B(pi03), .O(n410));
  andx g0312(.A(n2398), .B(n2461), .O(n411));
  andx g0313(.A(n225), .B(n2552), .O(n412));
  andx g0314(.A(n2668), .B(pi05), .O(n413));
  andx g0315(.A(n1126), .B(n2426), .O(n414));
  andx g0316(.A(n1083), .B(pi00), .O(n415));
  andx g0317(.A(n1125), .B(n2503), .O(n416));
  andx g0318(.A(n1127), .B(pi04), .O(n417));
  andx g0319(.A(pi03), .B(n2357), .O(n418));
  andx g0320(.A(n2398), .B(n2462), .O(n419));
  andx g0321(.A(n1130), .B(n1129), .O(n420));
  andx g0322(.A(n1132), .B(n1131), .O(n421));
  andx g0323(.A(n1128), .B(n2747), .O(n422));
  andx g0324(.A(n230), .B(pi06), .O(n423));
  andx g0325(.A(pi02), .B(n2461), .O(n424));
  andx g0326(.A(n2392), .B(pi03), .O(n425));
  andx g0327(.A(n2372), .B(n2463), .O(n426));
  andx g0328(.A(n2394), .B(pi03), .O(n427));
  andx g0329(.A(n237), .B(n2551), .O(n428));
  andx g0330(.A(n236), .B(pi05), .O(n429));
  andx g0331(.A(n2484), .B(n2358), .O(n430));
  andx g0332(.A(pi03), .B(n2383), .O(n431));
  andx g0333(.A(n2395), .B(n2462), .O(n432));
  andx g0334(.A(n2397), .B(pi03), .O(n433));
  andx g0335(.A(n235), .B(n2551), .O(n434));
  andx g0336(.A(n234), .B(pi05), .O(n435));
  andx g0337(.A(n1133), .B(n2426), .O(n436));
  andx g0338(.A(n1134), .B(pi00), .O(n437));
  andx g0339(.A(n2483), .B(n2330), .O(n438));
  andx g0340(.A(pi03), .B(n183), .O(n439));
  andx g0341(.A(pi01), .B(n2463), .O(n440));
  andx g0342(.A(pi03), .B(n2727), .O(n441));
  andx g0343(.A(n1136), .B(n2552), .O(n442));
  andx g0344(.A(n233), .B(pi05), .O(n443));
  andx g0345(.A(n2668), .B(pi05), .O(n444));
  andx g0346(.A(n2670), .B(n2552), .O(n445));
  andx g0347(.A(n1137), .B(n2426), .O(n446));
  andx g0348(.A(n1138), .B(pi00), .O(n447));
  andx g0349(.A(n1135), .B(n2503), .O(n448));
  andx g0350(.A(n1139), .B(pi04), .O(n449));
  andx g0351(.A(pi01), .B(n2462), .O(n450));
  andx g0352(.A(pi03), .B(n2355), .O(n451));
  andx g0353(.A(n1142), .B(n1141), .O(n452));
  andx g0354(.A(n232), .B(n2505), .O(n453));
  andx g0355(.A(n1084), .B(pi04), .O(n454));
  andx g0356(.A(n1140), .B(n2747), .O(n455));
  andx g0357(.A(n1143), .B(pi06), .O(n456));
  andx g0358(.A(n241), .B(pi05), .O(n457));
  andx g0359(.A(n240), .B(n2552), .O(n458));
  andx g0360(.A(n1085), .B(n2425), .O(n459));
  andx g0361(.A(n1144), .B(pi00), .O(n460));
  andx g0362(.A(n1086), .B(n2553), .O(n461));
  andx g0363(.A(n2601), .B(pi05), .O(n462));
  andx g0364(.A(n2369), .B(pi03), .O(n463));
  andx g0365(.A(n207), .B(n2464), .O(n464));
  andx g0366(.A(pi03), .B(n2359), .O(n465));
  andx g0367(.A(n2483), .B(n2760), .O(n466));
  andx g0368(.A(n1147), .B(n2553), .O(n467));
  andx g0369(.A(n239), .B(pi05), .O(n468));
  andx g0370(.A(n1146), .B(n2425), .O(n469));
  andx g0371(.A(n1148), .B(pi00), .O(n470));
  andx g0372(.A(n1145), .B(n2503), .O(n471));
  andx g0373(.A(n1149), .B(pi04), .O(n472));
  andx g0374(.A(n1152), .B(n1151), .O(n473));
  andx g0375(.A(pi03), .B(n2387), .O(n474));
  andx g0376(.A(n2377), .B(n2463), .O(n475));
  andx g0377(.A(n1154), .B(n1153), .O(n476));
  andx g0378(.A(n1156), .B(n1155), .O(n477));
  andx g0379(.A(n1150), .B(n2363), .O(n478));
  andx g0380(.A(n242), .B(pi06), .O(n479));
  andx g0381(.A(n2670), .B(n2553), .O(n480));
  andx g0382(.A(n245), .B(pi05), .O(n481));
  andx g0383(.A(pi05), .B(n2674), .O(n482));
  andx g0384(.A(n2667), .B(n2554), .O(n483));
  andx g0385(.A(n1157), .B(n2425), .O(n484));
  andx g0386(.A(n1158), .B(pi00), .O(n485));
  andx g0387(.A(n2659), .B(n2553), .O(n486));
  andx g0388(.A(n209), .B(pi05), .O(n487));
  andx g0389(.A(pi02), .B(n2464), .O(n488));
  andx g0390(.A(pi03), .B(n2370), .O(n489));
  andx g0391(.A(n2465), .B(n2358), .O(n490));
  andx g0392(.A(n2339), .B(pi03), .O(n491));
  andx g0393(.A(n1161), .B(n2554), .O(n492));
  andx g0394(.A(n1162), .B(pi05), .O(n493));
  andx g0395(.A(n1160), .B(n2425), .O(n494));
  andx g0396(.A(n1163), .B(pi00), .O(n495));
  andx g0397(.A(n1159), .B(n2523), .O(n496));
  andx g0398(.A(n1164), .B(pi04), .O(n497));
  andx g0399(.A(n1167), .B(n1166), .O(n498));
  andx g0400(.A(pi01), .B(n2463), .O(n499));
  andx g0401(.A(n2699), .B(pi03), .O(n500));
  andx g0402(.A(n1169), .B(n1168), .O(n501));
  andx g0403(.A(n1171), .B(n1170), .O(n502));
  andx g0404(.A(n1165), .B(n2352), .O(n503));
  andx g0405(.A(n246), .B(pi06), .O(n504));
  andx g0406(.A(n2658), .B(n2554), .O(n505));
  andx g0407(.A(n2652), .B(pi05), .O(n506));
  andx g0408(.A(pi03), .B(n2348), .O(n507));
  andx g0409(.A(n2338), .B(n2465), .O(n508));
  andx g0410(.A(pi03), .B(n2356), .O(n509));
  andx g0411(.A(n2385), .B(n2464), .O(n510));
  andx g0412(.A(n1173), .B(n2555), .O(n511));
  andx g0413(.A(n1174), .B(pi05), .O(n512));
  andx g0414(.A(n1172), .B(n2424), .O(n513));
  andx g0415(.A(n1175), .B(pi00), .O(n514));
  andx g0416(.A(n2461), .B(n2357), .O(n515));
  andx g0417(.A(pi03), .B(n2385), .O(n516));
  andx g0418(.A(n191), .B(n2555), .O(n517));
  andx g0419(.A(n249), .B(pi05), .O(n518));
  andx g0420(.A(pi05), .B(n186), .O(n519));
  andx g0421(.A(n2655), .B(n2555), .O(n520));
  andx g0422(.A(n1177), .B(n2424), .O(n521));
  andx g0423(.A(n1178), .B(pi00), .O(n522));
  andx g0424(.A(n1176), .B(n2504), .O(n523));
  andx g0425(.A(n1179), .B(pi04), .O(n524));
  andx g0426(.A(n2483), .B(n2356), .O(n525));
  andx g0427(.A(n2378), .B(pi03), .O(n526));
  andx g0428(.A(n1182), .B(n1181), .O(n527));
  andx g0429(.A(n1184), .B(n1183), .O(n528));
  andx g0430(.A(n1186), .B(n1185), .O(n529));
  andx g0431(.A(n1180), .B(n2747), .O(n530));
  andx g0432(.A(n250), .B(pi06), .O(n531));
  andx g0433(.A(n1187), .B(n1188), .O(n532));
  andx g0434(.A(n2339), .B(n2555), .O(n533));
  andx g0435(.A(n254), .B(pi05), .O(n534));
  andx g0436(.A(n255), .B(n2424), .O(n535));
  andx g0437(.A(n1189), .B(pi00), .O(n536));
  orx  g0438(.A(n2598), .B(n2350), .O(n537));
  andx g0439(.A(n1192), .B(n1191), .O(n538));
  andx g0440(.A(n1194), .B(n1193), .O(n539));
  andx g0441(.A(n1196), .B(n1195), .O(n540));
  andx g0442(.A(n217), .B(pi06), .O(n541));
  andx g0443(.A(n540), .B(n2352), .O(n542));
  andx g0444(.A(n1197), .B(n2556), .O(n543));
  andx g0445(.A(n252), .B(pi05), .O(n544));
  andx g0446(.A(n253), .B(n2424), .O(n545));
  andx g0447(.A(n1198), .B(pi00), .O(n546));
  andx g0448(.A(n1190), .B(n2509), .O(n547));
  andx g0449(.A(n1199), .B(pi04), .O(n548));
  andx g0450(.A(pi01), .B(pi03), .O(n549));
  andx g0451(.A(n2397), .B(n2465), .O(n550));
  andx g0452(.A(n221), .B(n2751), .O(n551));
  andx g0453(.A(n1200), .B(pi04), .O(n552));
  orx  g0454(.A(n2338), .B(n2660), .O(n553));
  andx g0455(.A(pi04), .B(n203), .O(n554));
  andx g0456(.A(n2661), .B(n2504), .O(n555));
  andx g0457(.A(n1201), .B(n2423), .O(n556));
  andx g0458(.A(n1202), .B(pi00), .O(n557));
  andx g0459(.A(n2654), .B(pi04), .O(n558));
  andx g0460(.A(n2649), .B(n2504), .O(n559));
  andx g0461(.A(n2757), .B(n2360), .O(n560));
  andx g0462(.A(n2373), .B(pi03), .O(n561));
  andx g0463(.A(n209), .B(pi04), .O(n562));
  andx g0464(.A(n1205), .B(n2506), .O(n563));
  andx g0465(.A(n1204), .B(n2423), .O(n564));
  andx g0466(.A(n1206), .B(pi00), .O(n565));
  andx g0467(.A(n1203), .B(n2556), .O(n566));
  andx g0468(.A(n1207), .B(pi05), .O(n567));
  andx g0469(.A(n1210), .B(n1209), .O(n568));
  andx g0470(.A(n228), .B(pi04), .O(n569));
  andx g0471(.A(n175), .B(n2505), .O(n570));
  andx g0472(.A(n1212), .B(n1211), .O(n571));
  andx g0473(.A(n1208), .B(n2331), .O(n572));
  andx g0474(.A(n258), .B(pi06), .O(n573));
  andx g0475(.A(pi03), .B(n2764), .O(n574));
  andx g0476(.A(n2338), .B(n2464), .O(n575));
  andx g0477(.A(pi05), .B(n201), .O(n576));
  andx g0478(.A(n1213), .B(n2556), .O(n577));
  andx g0479(.A(n186), .B(n2556), .O(n578));
  andx g0480(.A(n226), .B(pi05), .O(n579));
  andx g0481(.A(n1214), .B(n2423), .O(n580));
  andx g0482(.A(n1215), .B(pi00), .O(n581));
  andx g0483(.A(n2483), .B(n2354), .O(n582));
  andx g0484(.A(n2368), .B(pi03), .O(n583));
  orx  g0485(.A(n2609), .B(n2384), .O(n584));
  andx g0486(.A(n2610), .B(n2557), .O(n585));
  andx g0487(.A(n262), .B(pi05), .O(n586));
  andx g0488(.A(pi03), .B(n2358), .O(n587));
  andx g0489(.A(n2387), .B(n2466), .O(n588));
  andx g0490(.A(n221), .B(n2557), .O(n589));
  andx g0491(.A(n261), .B(pi05), .O(n590));
  andx g0492(.A(n1217), .B(n2423), .O(n591));
  andx g0493(.A(n1218), .B(pi00), .O(n592));
  andx g0494(.A(n1216), .B(n2505), .O(n593));
  andx g0495(.A(n1219), .B(pi04), .O(n594));
  andx g0496(.A(n1222), .B(n1221), .O(n595));
  orx  g0497(.A(pi05), .B(n202), .O(n596));
  andx g0498(.A(n2711), .B(n2422), .O(n597));
  andx g0499(.A(n2628), .B(pi00), .O(n598));
  andx g0500(.A(n260), .B(n2507), .O(n599));
  andx g0501(.A(n1223), .B(pi04), .O(n600));
  andx g0502(.A(n1220), .B(n2351), .O(n601));
  andx g0503(.A(n1224), .B(pi06), .O(n602));
  andx g0504(.A(n2482), .B(n2360), .O(n603));
  andx g0505(.A(n2369), .B(pi03), .O(n604));
  andx g0506(.A(n244), .B(n2557), .O(n605));
  andx g0507(.A(n1225), .B(pi05), .O(n606));
  andx g0508(.A(n239), .B(pi05), .O(n607));
  andx g0509(.A(n2631), .B(n2557), .O(n608));
  andx g0510(.A(n1226), .B(n2415), .O(n609));
  andx g0511(.A(n1227), .B(pi00), .O(n610));
  andx g0512(.A(n2647), .B(n2558), .O(n611));
  andx g0513(.A(n240), .B(pi05), .O(n612));
  andx g0514(.A(pi01), .B(pi03), .O(n613));
  andx g0515(.A(n2393), .B(n2465), .O(n614));
  andx g0516(.A(n2368), .B(pi05), .O(n615));
  andx g0517(.A(n1230), .B(n2558), .O(n616));
  andx g0518(.A(n1229), .B(n2422), .O(n617));
  andx g0519(.A(n1231), .B(pi00), .O(n618));
  andx g0520(.A(n1228), .B(n2508), .O(n619));
  andx g0521(.A(n1232), .B(pi04), .O(n620));
  andx g0522(.A(n1235), .B(n1234), .O(n621));
  andx g0523(.A(n1237), .B(n1236), .O(n622));
  andx g0524(.A(n1233), .B(n2349), .O(n623));
  andx g0525(.A(n264), .B(pi06), .O(n624));
  andx g0526(.A(n208), .B(n2558), .O(n625));
  andx g0527(.A(pi05), .B(n199), .O(n626));
  andx g0528(.A(n172), .B(pi05), .O(n627));
  andx g0529(.A(n2729), .B(n2558), .O(n628));
  andx g0530(.A(n1238), .B(n2422), .O(n629));
  andx g0531(.A(n1239), .B(pi00), .O(n630));
  andx g0532(.A(n2347), .B(n2466), .O(n631));
  andx g0533(.A(n2369), .B(pi03), .O(n632));
  andx g0534(.A(n175), .B(pi05), .O(n633));
  andx g0535(.A(n1241), .B(n2559), .O(n634));
  andx g0536(.A(pi01), .B(n2465), .O(n635));
  andx g0537(.A(n2392), .B(pi03), .O(n636));
  andx g0538(.A(pi05), .B(n185), .O(n637));
  andx g0539(.A(n269), .B(n2559), .O(n638));
  andx g0540(.A(n1242), .B(n2421), .O(n639));
  andx g0541(.A(n1243), .B(pi00), .O(n640));
  andx g0542(.A(n1240), .B(n2505), .O(n641));
  andx g0543(.A(n1244), .B(pi04), .O(n642));
  andx g0544(.A(pi03), .B(n2361), .O(n643));
  andx g0545(.A(n2366), .B(n2467), .O(n644));
  orx  g0546(.A(n2397), .B(n2485), .O(n645));
  andx g0547(.A(n1247), .B(n1246), .O(n646));
  andx g0548(.A(n2384), .B(n2466), .O(n647));
  andx g0549(.A(n2377), .B(pi03), .O(n648));
  orx  g0550(.A(pi05), .B(n191), .O(n649));
  orx  g0551(.A(pi05), .B(n2625), .O(n650));
  andx g0552(.A(n2702), .B(n2421), .O(n651));
  andx g0553(.A(n2694), .B(pi00), .O(n652));
  andx g0554(.A(n268), .B(n2508), .O(n653));
  andx g0555(.A(n1248), .B(pi04), .O(n654));
  andx g0556(.A(n1245), .B(n2362), .O(n655));
  andx g0557(.A(n1249), .B(pi06), .O(n656));
  andx g0558(.A(pi03), .B(n2356), .O(n657));
  andx g0559(.A(n2348), .B(n2467), .O(n658));
  andx g0560(.A(n172), .B(n2559), .O(n659));
  andx g0561(.A(n1250), .B(pi05), .O(n660));
  andx g0562(.A(n2372), .B(n2466), .O(n661));
  andx g0563(.A(n2398), .B(pi03), .O(n662));
  andx g0564(.A(n2699), .B(n2559), .O(n663));
  andx g0565(.A(n272), .B(pi05), .O(n664));
  andx g0566(.A(n1251), .B(n2421), .O(n665));
  andx g0567(.A(n1252), .B(pi00), .O(n666));
  andx g0568(.A(n2600), .B(pi05), .O(n667));
  andx g0569(.A(n176), .B(n2560), .O(n668));
  andx g0570(.A(n236), .B(n2560), .O(n669));
  andx g0571(.A(n2630), .B(pi05), .O(n670));
  andx g0572(.A(n1254), .B(n2421), .O(n671));
  andx g0573(.A(n1255), .B(pi00), .O(n672));
  andx g0574(.A(n1253), .B(n2522), .O(n673));
  andx g0575(.A(n1256), .B(pi04), .O(n674));
  andx g0576(.A(n1259), .B(n1258), .O(n675));
  orx  g0577(.A(pi05), .B(n197), .O(n676));
  andx g0578(.A(n2607), .B(n2420), .O(n677));
  andx g0579(.A(n2685), .B(pi00), .O(n678));
  andx g0580(.A(n271), .B(n2751), .O(n679));
  andx g0581(.A(n1260), .B(pi04), .O(n680));
  andx g0582(.A(n1257), .B(n2335), .O(n681));
  andx g0583(.A(n1261), .B(pi06), .O(n682));
  orx  g0584(.A(n2457), .B(n2760), .O(n683));
  andx g0585(.A(n2645), .B(pi05), .O(n684));
  andx g0586(.A(n2623), .B(n2560), .O(n685));
  andx g0587(.A(n2339), .B(n2467), .O(n686));
  andx g0588(.A(pi03), .B(n2384), .O(n687));
  andx g0589(.A(pi02), .B(pi03), .O(n688));
  andx g0590(.A(n2373), .B(n2468), .O(n689));
  andx g0591(.A(n277), .B(n2560), .O(n690));
  andx g0592(.A(n276), .B(pi05), .O(n691));
  andx g0593(.A(n1262), .B(n2420), .O(n692));
  andx g0594(.A(n1263), .B(pi00), .O(n693));
  andx g0595(.A(n1112), .B(n2561), .O(n694));
  andx g0596(.A(n236), .B(pi05), .O(n695));
  andx g0597(.A(n2658), .B(n2561), .O(n696));
  andx g0598(.A(pi05), .B(n191), .O(n697));
  andx g0599(.A(n1265), .B(n2420), .O(n698));
  andx g0600(.A(n1266), .B(pi00), .O(n699));
  andx g0601(.A(n1264), .B(n2508), .O(n700));
  andx g0602(.A(n1267), .B(pi04), .O(n701));
  andx g0603(.A(pi01), .B(pi03), .O(n702));
  andx g0604(.A(n2387), .B(n2471), .O(n703));
  andx g0605(.A(n1270), .B(n1269), .O(n704));
  andx g0606(.A(n2639), .B(pi00), .O(n705));
  andx g0607(.A(n2711), .B(n2420), .O(n706));
  andx g0608(.A(n275), .B(n2506), .O(n707));
  andx g0609(.A(n1271), .B(pi04), .O(n708));
  andx g0610(.A(n1268), .B(n2353), .O(n709));
  andx g0611(.A(n1272), .B(pi06), .O(n710));
  orx  g0612(.A(n2377), .B(n2626), .O(n711));
  andx g0613(.A(n1082), .B(pi05), .O(n712));
  andx g0614(.A(n2627), .B(n2561), .O(n713));
  andx g0615(.A(pi03), .B(n2346), .O(n714));
  andx g0616(.A(n2395), .B(n2467), .O(n715));
  andx g0617(.A(n1274), .B(n2561), .O(n716));
  andx g0618(.A(n2611), .B(pi05), .O(n717));
  andx g0619(.A(n1273), .B(n2419), .O(n718));
  andx g0620(.A(n1275), .B(pi00), .O(n719));
  andx g0621(.A(n212), .B(pi05), .O(n720));
  andx g0622(.A(n229), .B(n2562), .O(n721));
  andx g0623(.A(n2652), .B(pi05), .O(n722));
  andx g0624(.A(n199), .B(n2562), .O(n723));
  andx g0625(.A(n1277), .B(n2419), .O(n724));
  andx g0626(.A(n1278), .B(pi00), .O(n725));
  andx g0627(.A(n1276), .B(n2506), .O(n726));
  andx g0628(.A(n1279), .B(pi04), .O(n727));
  andx g0629(.A(pi03), .B(n2330), .O(n728));
  andx g0630(.A(n2397), .B(n2468), .O(n729));
  andx g0631(.A(n2482), .B(n2360), .O(n730));
  andx g0632(.A(n2378), .B(pi03), .O(n731));
  andx g0633(.A(n1282), .B(n1281), .O(n732));
  andx g0634(.A(n2702), .B(pi00), .O(n733));
  andx g0635(.A(n2711), .B(n2419), .O(n734));
  andx g0636(.A(n281), .B(n2510), .O(n735));
  andx g0637(.A(n1283), .B(pi04), .O(n736));
  andx g0638(.A(n1280), .B(n2747), .O(n737));
  andx g0639(.A(n1284), .B(pi06), .O(n738));
  andx g0640(.A(n2600), .B(pi05), .O(n739));
  andx g0641(.A(n2624), .B(n2562), .O(n740));
  andx g0642(.A(n2652), .B(pi05), .O(n741));
  andx g0643(.A(n2671), .B(n2562), .O(n742));
  andx g0644(.A(n1285), .B(n2419), .O(n743));
  andx g0645(.A(n1286), .B(pi00), .O(n744));
  andx g0646(.A(pi03), .B(n2361), .O(n745));
  andx g0647(.A(n2368), .B(n2468), .O(n746));
  andx g0648(.A(n2665), .B(n2563), .O(n747));
  andx g0649(.A(n284), .B(pi05), .O(n748));
  andx g0650(.A(pi01), .B(n2469), .O(n749));
  andx g0651(.A(pi03), .B(n2383), .O(n750));
  andx g0652(.A(n1288), .B(n2418), .O(n751));
  andx g0653(.A(n1088), .B(pi00), .O(n752));
  andx g0654(.A(n1287), .B(n2506), .O(n753));
  andx g0655(.A(n1289), .B(pi04), .O(n754));
  andx g0656(.A(n1292), .B(n1291), .O(n755));
  andx g0657(.A(n1294), .B(n1293), .O(n756));
  andx g0658(.A(n1296), .B(n1295), .O(n757));
  andx g0659(.A(n1290), .B(n2747), .O(n758));
  andx g0660(.A(n285), .B(pi06), .O(n759));
  andx g0661(.A(pi05), .B(n2666), .O(n760));
  andx g0662(.A(n2621), .B(n2563), .O(n761));
  andx g0663(.A(pi05), .B(n2727), .O(n762));
  andx g0664(.A(n2629), .B(n2563), .O(n763));
  andx g0665(.A(n1297), .B(n2418), .O(n764));
  andx g0666(.A(n1298), .B(pi00), .O(n765));
  andx g0667(.A(pi01), .B(n2468), .O(n766));
  andx g0668(.A(n2338), .B(pi03), .O(n767));
  andx g0669(.A(n1230), .B(pi05), .O(n768));
  andx g0670(.A(n288), .B(n2563), .O(n769));
  andx g0671(.A(n165), .B(n2564), .O(n770));
  andx g0672(.A(n2629), .B(pi05), .O(n771));
  andx g0673(.A(n1300), .B(n2418), .O(n772));
  andx g0674(.A(n1301), .B(pi00), .O(n773));
  andx g0675(.A(n1299), .B(n2507), .O(n774));
  andx g0676(.A(n1302), .B(pi04), .O(n775));
  orx  g0677(.A(pi05), .B(n2634), .O(n776));
  andx g0678(.A(n287), .B(n2418), .O(n777));
  andx g0679(.A(n2684), .B(pi00), .O(n778));
  andx g0680(.A(n2731), .B(pi04), .O(n779));
  andx g0681(.A(n1304), .B(n2510), .O(n780));
  andx g0682(.A(n1303), .B(n2349), .O(n781));
  andx g0683(.A(n1305), .B(pi06), .O(n782));
  andx g0684(.A(n2675), .B(pi05), .O(n783));
  andx g0685(.A(n207), .B(n2564), .O(n784));
  andx g0686(.A(n274), .B(n2564), .O(n785));
  andx g0687(.A(n291), .B(pi05), .O(n786));
  andx g0688(.A(n1306), .B(n2417), .O(n787));
  andx g0689(.A(n1307), .B(pi00), .O(n788));
  andx g0690(.A(n215), .B(n2564), .O(n789));
  andx g0691(.A(n2600), .B(pi05), .O(n790));
  andx g0692(.A(n2584), .B(n2760), .O(n791));
  andx g0693(.A(pi05), .B(n201), .O(n792));
  andx g0694(.A(n1309), .B(n2428), .O(n793));
  andx g0695(.A(n1310), .B(pi00), .O(n794));
  andx g0696(.A(n1308), .B(n2507), .O(n795));
  andx g0697(.A(n1311), .B(pi04), .O(n796));
  andx g0698(.A(n1314), .B(n1313), .O(n797));
  andx g0699(.A(n1316), .B(n1315), .O(n798));
  andx g0700(.A(n2607), .B(pi00), .O(n799));
  andx g0701(.A(n2617), .B(n2417), .O(n800));
  andx g0702(.A(n290), .B(n2507), .O(n801));
  andx g0703(.A(n1317), .B(pi04), .O(n802));
  andx g0704(.A(n1312), .B(n2352), .O(n803));
  andx g0705(.A(n1318), .B(pi06), .O(n804));
  andx g0706(.A(pi01), .B(n2469), .O(n805));
  andx g0707(.A(n2369), .B(pi03), .O(n806));
  andx g0708(.A(n2610), .B(pi05), .O(n807));
  andx g0709(.A(n294), .B(n2562), .O(n808));
  andx g0710(.A(n2398), .B(pi05), .O(n809));
  andx g0711(.A(n2632), .B(n2554), .O(n810));
  andx g0712(.A(n1319), .B(n2417), .O(n811));
  andx g0713(.A(n1320), .B(pi00), .O(n812));
  andx g0714(.A(n163), .B(n2553), .O(n813));
  andx g0715(.A(n274), .B(pi05), .O(n814));
  andx g0716(.A(n198), .B(n2565), .O(n815));
  andx g0717(.A(n269), .B(pi05), .O(n816));
  andx g0718(.A(n1322), .B(n2417), .O(n817));
  andx g0719(.A(n1323), .B(pi00), .O(n818));
  andx g0720(.A(n1321), .B(n2511), .O(n819));
  andx g0721(.A(n1324), .B(pi04), .O(n820));
  andx g0722(.A(n1327), .B(n1326), .O(n821));
  andx g0723(.A(n1329), .B(n1328), .O(n822));
  andx g0724(.A(n2731), .B(pi00), .O(n823));
  andx g0725(.A(n2617), .B(n2416), .O(n824));
  andx g0726(.A(n293), .B(n2508), .O(n825));
  andx g0727(.A(n1330), .B(pi04), .O(n826));
  andx g0728(.A(n1325), .B(n2336), .O(n827));
  andx g0729(.A(n1331), .B(pi06), .O(n828));
  andx g0730(.A(pi02), .B(n2469), .O(n829));
  andx g0731(.A(pi03), .B(n2359), .O(n830));
  andx g0732(.A(n1200), .B(pi04), .O(n831));
  andx g0733(.A(n211), .B(n2516), .O(n832));
  andx g0734(.A(pi04), .B(pi02), .O(n833));
  andx g0735(.A(n219), .B(n2511), .O(n834));
  andx g0736(.A(n1332), .B(n2416), .O(n835));
  andx g0737(.A(n1333), .B(pi00), .O(n836));
  andx g0738(.A(n2662), .B(n2509), .O(n837));
  andx g0739(.A(n1089), .B(pi04), .O(n838));
  andx g0740(.A(n1335), .B(n2416), .O(n839));
  andx g0741(.A(n296), .B(pi00), .O(n840));
  andx g0742(.A(n1334), .B(n2565), .O(n841));
  andx g0743(.A(n1336), .B(pi05), .O(n842));
  andx g0744(.A(n1339), .B(n1338), .O(n843));
  orx  g0745(.A(n2606), .B(n2530), .O(n844));
  andx g0746(.A(n1341), .B(n1340), .O(n845));
  andx g0747(.A(n1337), .B(n2335), .O(n846));
  andx g0748(.A(n297), .B(pi06), .O(n847));
  andx g0749(.A(n2604), .B(n2416), .O(n848));
  andx g0750(.A(n2623), .B(pi00), .O(n849));
  andx g0751(.A(n2657), .B(n2415), .O(n850));
  andx g0752(.A(n1091), .B(pi00), .O(n851));
  andx g0753(.A(n1342), .B(n2509), .O(n852));
  andx g0754(.A(n1343), .B(pi04), .O(n853));
  andx g0755(.A(n2640), .B(n2415), .O(n854));
  andx g0756(.A(n1250), .B(pi00), .O(n855));
  orx  g0757(.A(n2668), .B(n2383), .O(n856));
  andx g0758(.A(n2634), .B(pi00), .O(n857));
  andx g0759(.A(n2669), .B(n2415), .O(n858));
  andx g0760(.A(n1345), .B(n2512), .O(n859));
  andx g0761(.A(n1346), .B(pi04), .O(n860));
  andx g0762(.A(n1344), .B(n2565), .O(n861));
  andx g0763(.A(n1347), .B(pi05), .O(n862));
  andx g0764(.A(pi02), .B(n2470), .O(n863));
  andx g0765(.A(n2368), .B(pi03), .O(n864));
  andx g0766(.A(n1350), .B(n1349), .O(n865));
  andx g0767(.A(n1352), .B(n1351), .O(n866));
  andx g0768(.A(n1354), .B(n1353), .O(n867));
  andx g0769(.A(n1348), .B(n2350), .O(n868));
  andx g0770(.A(n300), .B(pi06), .O(n869));
  andx g0771(.A(pi04), .B(n2672), .O(n870));
  andx g0772(.A(n2621), .B(n2509), .O(n871));
  andx g0773(.A(n2682), .B(n2414), .O(n872));
  andx g0774(.A(n1355), .B(pi00), .O(n873));
  andx g0775(.A(n196), .B(n2510), .O(n874));
  andx g0776(.A(n262), .B(pi04), .O(n875));
  andx g0777(.A(n2655), .B(n2513), .O(n876));
  andx g0778(.A(n2642), .B(pi04), .O(n877));
  andx g0779(.A(n1357), .B(n2414), .O(n878));
  andx g0780(.A(n1358), .B(pi00), .O(n879));
  andx g0781(.A(n1356), .B(n2565), .O(n880));
  andx g0782(.A(n1359), .B(pi05), .O(n881));
  andx g0783(.A(n1362), .B(n1361), .O(n882));
  andx g0784(.A(n1364), .B(n1363), .O(n883));
  andx g0785(.A(n1360), .B(n2351), .O(n884));
  andx g0786(.A(n303), .B(pi06), .O(n885));
  andx g0787(.A(pi05), .B(n205), .O(n886));
  andx g0788(.A(n2619), .B(n2566), .O(n887));
  andx g0789(.A(n1273), .B(pi00), .O(n888));
  andx g0790(.A(n1365), .B(n2414), .O(n889));
  andx g0791(.A(n2339), .B(n2566), .O(n890));
  andx g0792(.A(pi05), .B(n193), .O(n891));
  andx g0793(.A(n1367), .B(n2414), .O(n892));
  andx g0794(.A(n306), .B(pi00), .O(n893));
  andx g0795(.A(n1366), .B(n2515), .O(n894));
  andx g0796(.A(n1368), .B(pi04), .O(n895));
  andx g0797(.A(n1371), .B(n1370), .O(n896));
  andx g0798(.A(n2711), .B(n2765), .O(n897));
  andx g0799(.A(n2617), .B(pi00), .O(n898));
  andx g0800(.A(n305), .B(n2510), .O(n899));
  andx g0801(.A(n1372), .B(pi04), .O(n900));
  andx g0802(.A(n1369), .B(n2353), .O(n901));
  andx g0803(.A(n1373), .B(pi06), .O(n902));
  andx g0804(.A(n2653), .B(pi05), .O(n903));
  andx g0805(.A(n2624), .B(n2566), .O(n904));
  andx g0806(.A(n2623), .B(pi05), .O(n905));
  andx g0807(.A(n2622), .B(n2566), .O(n906));
  andx g0808(.A(n1374), .B(n2765), .O(n907));
  andx g0809(.A(n1375), .B(pi00), .O(n908));
  andx g0810(.A(pi05), .B(n2355), .O(n909));
  andx g0811(.A(n276), .B(n2567), .O(n910));
  andx g0812(.A(n1218), .B(n2437), .O(n911));
  andx g0813(.A(n1377), .B(pi00), .O(n912));
  andx g0814(.A(n1376), .B(n2514), .O(n913));
  andx g0815(.A(n1378), .B(pi04), .O(n914));
  andx g0816(.A(n2711), .B(pi00), .O(n915));
  andx g0817(.A(n2685), .B(n2438), .O(n916));
  andx g0818(.A(n2694), .B(pi00), .O(n917));
  andx g0819(.A(n2684), .B(n2413), .O(n918));
  andx g0820(.A(n1380), .B(n2511), .O(n919));
  andx g0821(.A(n1381), .B(pi04), .O(n920));
  andx g0822(.A(n1379), .B(n2363), .O(n921));
  andx g0823(.A(n1382), .B(pi06), .O(n922));
  andx g0824(.A(pi03), .B(n2764), .O(n923));
  andx g0825(.A(n2377), .B(n2469), .O(n924));
  andx g0826(.A(n192), .B(n2567), .O(n925));
  andx g0827(.A(n1383), .B(pi05), .O(n926));
  andx g0828(.A(n310), .B(n2413), .O(n927));
  andx g0829(.A(n1384), .B(pi00), .O(n928));
  andx g0830(.A(n1225), .B(n2567), .O(n929));
  andx g0831(.A(n299), .B(pi05), .O(n930));
  andx g0832(.A(n2641), .B(pi05), .O(n931));
  andx g0833(.A(n2616), .B(n2567), .O(n932));
  andx g0834(.A(n1386), .B(n2413), .O(n933));
  andx g0835(.A(n1387), .B(pi00), .O(n934));
  andx g0836(.A(n1385), .B(n2511), .O(n935));
  andx g0837(.A(n1388), .B(pi04), .O(n936));
  andx g0838(.A(n1391), .B(n1390), .O(n937));
  andx g0839(.A(n309), .B(n2514), .O(n938));
  andx g0840(.A(n1095), .B(pi04), .O(n939));
  andx g0841(.A(n1389), .B(n2363), .O(n940));
  andx g0842(.A(n1392), .B(pi06), .O(n941));
  andx g0843(.A(n190), .B(n2568), .O(n942));
  andx g0844(.A(pi05), .B(n192), .O(n943));
  andx g0845(.A(n2584), .B(n2354), .O(n944));
  andx g0846(.A(pi05), .B(n2370), .O(n945));
  andx g0847(.A(n2699), .B(n2470), .O(n946));
  andx g0848(.A(n1394), .B(pi03), .O(n947));
  andx g0849(.A(n1393), .B(n2413), .O(n948));
  andx g0850(.A(n1395), .B(pi00), .O(n949));
  andx g0851(.A(pi01), .B(n2568), .O(n950));
  andx g0852(.A(n274), .B(pi05), .O(n951));
  andx g0853(.A(n2651), .B(n2568), .O(n952));
  andx g0854(.A(pi05), .B(n205), .O(n953));
  andx g0855(.A(n1397), .B(n2412), .O(n954));
  andx g0856(.A(n1398), .B(pi00), .O(n955));
  andx g0857(.A(n1396), .B(n2512), .O(n956));
  andx g0858(.A(n1399), .B(pi04), .O(n957));
  andx g0859(.A(n1402), .B(n1401), .O(n958));
  andx g0860(.A(n1404), .B(n1403), .O(n959));
  andx g0861(.A(n1406), .B(n1405), .O(n960));
  andx g0862(.A(n1400), .B(n2353), .O(n961));
  andx g0863(.A(n312), .B(pi06), .O(n962));
  andx g0864(.A(pi01), .B(pi03), .O(n963));
  andx g0865(.A(n2347), .B(n2470), .O(n964));
  andx g0866(.A(n201), .B(n2568), .O(n965));
  andx g0867(.A(n315), .B(pi05), .O(n966));
  andx g0868(.A(n1173), .B(n2569), .O(n967));
  andx g0869(.A(n2669), .B(pi05), .O(n968));
  andx g0870(.A(n1407), .B(n2412), .O(n969));
  andx g0871(.A(n1408), .B(pi00), .O(n970));
  andx g0872(.A(n1082), .B(n2569), .O(n971));
  andx g0873(.A(n2626), .B(pi05), .O(n972));
  andx g0874(.A(n2348), .B(n2470), .O(n973));
  andx g0875(.A(pi03), .B(n2386), .O(n974));
  andx g0876(.A(n2584), .B(n2760), .O(n975));
  andx g0877(.A(n1411), .B(pi05), .O(n976));
  andx g0878(.A(n1410), .B(n2412), .O(n977));
  andx g0879(.A(n1412), .B(pi00), .O(n978));
  andx g0880(.A(n1409), .B(n2512), .O(n979));
  andx g0881(.A(n1413), .B(pi04), .O(n980));
  andx g0882(.A(n1416), .B(n1415), .O(n981));
  andx g0883(.A(n314), .B(n2514), .O(n982));
  andx g0884(.A(n1096), .B(pi04), .O(n983));
  andx g0885(.A(n1414), .B(n2349), .O(n984));
  andx g0886(.A(n1417), .B(pi06), .O(n985));
  andx g0887(.A(pi05), .B(n2605), .O(n986));
  andx g0888(.A(n2627), .B(n2570), .O(n987));
  andx g0889(.A(pi05), .B(n2385), .O(n988));
  andx g0890(.A(n184), .B(n2570), .O(n989));
  andx g0891(.A(n1418), .B(n2411), .O(n990));
  andx g0892(.A(n1419), .B(pi00), .O(n991));
  andx g0893(.A(n237), .B(pi05), .O(n992));
  andx g0894(.A(n2615), .B(n2569), .O(n993));
  andx g0895(.A(n1229), .B(n2411), .O(n994));
  andx g0896(.A(n1421), .B(pi00), .O(n995));
  andx g0897(.A(n1420), .B(n2512), .O(n996));
  andx g0898(.A(n1422), .B(pi04), .O(n997));
  andx g0899(.A(n1425), .B(n1424), .O(n998));
  andx g0900(.A(n1427), .B(n1426), .O(n999));
  andx g0901(.A(n1429), .B(n1428), .O(n1000));
  andx g0902(.A(n1431), .B(n1430), .O(n1001));
  andx g0903(.A(n1423), .B(n2747), .O(n1002));
  andx g0904(.A(n317), .B(pi06), .O(n1003));
  andx g0905(.A(n2648), .B(pi05), .O(n1004));
  andx g0906(.A(n190), .B(n2570), .O(n1005));
  andx g0907(.A(pi05), .B(n2673), .O(n1006));
  andx g0908(.A(n205), .B(n2571), .O(n1007));
  andx g0909(.A(n1432), .B(n2411), .O(n1008));
  andx g0910(.A(n1433), .B(pi00), .O(n1009));
  andx g0911(.A(n2598), .B(pi05), .O(n1010));
  andx g0912(.A(n1411), .B(n2569), .O(n1011));
  andx g0913(.A(n217), .B(n2571), .O(n1012));
  andx g0914(.A(n2649), .B(pi05), .O(n1013));
  andx g0915(.A(n1435), .B(n2410), .O(n1014));
  andx g0916(.A(n1436), .B(pi00), .O(n1015));
  andx g0917(.A(n1434), .B(n2513), .O(n1016));
  andx g0918(.A(n1437), .B(pi04), .O(n1017));
  andx g0919(.A(n1440), .B(n1439), .O(n1018));
  andx g0920(.A(n1442), .B(n1441), .O(n1019));
  andx g0921(.A(n1444), .B(n1443), .O(n1020));
  andx g0922(.A(n1438), .B(n2350), .O(n1021));
  andx g0923(.A(n319), .B(pi06), .O(n1022));
  andx g0924(.A(n2372), .B(pi03), .O(n1023));
  andx g0925(.A(n2386), .B(n2471), .O(n1024));
  andx g0926(.A(n194), .B(n2515), .O(n1025));
  andx g0927(.A(n1445), .B(pi04), .O(n1026));
  andx g0928(.A(n2527), .B(n2357), .O(n1027));
  andx g0929(.A(pi04), .B(n186), .O(n1028));
  andx g0930(.A(n1446), .B(n2410), .O(n1029));
  andx g0931(.A(n1447), .B(pi00), .O(n1030));
  andx g0932(.A(n2646), .B(pi04), .O(n1031));
  andx g0933(.A(n2620), .B(n2513), .O(n1032));
  andx g0934(.A(n2655), .B(pi04), .O(n1033));
  andx g0935(.A(n187), .B(n2513), .O(n1034));
  andx g0936(.A(n1449), .B(n2412), .O(n1035));
  andx g0937(.A(n1450), .B(pi00), .O(n1036));
  andx g0938(.A(n1448), .B(n2571), .O(n1037));
  andx g0939(.A(n1451), .B(pi05), .O(n1038));
  andx g0940(.A(n1454), .B(n1453), .O(n1039));
  andx g0941(.A(n1456), .B(n1455), .O(n1040));
  andx g0942(.A(n1458), .B(n1457), .O(n1041));
  andx g0943(.A(n1452), .B(n2352), .O(n1042));
  andx g0944(.A(n321), .B(pi06), .O(n1043));
  andx g0945(.A(n1200), .B(n2515), .O(n1044));
  andx g0946(.A(n2625), .B(pi04), .O(n1045));
  andx g0947(.A(n2655), .B(pi04), .O(n1046));
  andx g0948(.A(n269), .B(n2514), .O(n1047));
  andx g0949(.A(n1459), .B(n2422), .O(n1048));
  andx g0950(.A(n1460), .B(pi00), .O(n1049));
  andx g0951(.A(n2658), .B(pi04), .O(n1050));
  andx g0952(.A(n2614), .B(n2515), .O(n1051));
  andx g0953(.A(n1097), .B(n2428), .O(n1052));
  andx g0954(.A(n1462), .B(pi00), .O(n1053));
  andx g0955(.A(n1461), .B(n2570), .O(n1054));
  andx g0956(.A(n1463), .B(pi05), .O(n1055));
  andx g0957(.A(n1466), .B(n1465), .O(n1056));
  andx g0958(.A(n1468), .B(n1467), .O(n1057));
  andx g0959(.A(n1470), .B(n1469), .O(n1058));
  andx g0960(.A(n1464), .B(n2363), .O(n1059));
  andx g0961(.A(n323), .B(pi06), .O(n1060));
  andx g0962(.A(pi05), .B(pi01), .O(n1061));
  andx g0963(.A(n2635), .B(n2572), .O(n1062));
  andx g0964(.A(n2654), .B(n2572), .O(n1063));
  andx g0965(.A(pi05), .B(n1081), .O(n1064));
  andx g0966(.A(n1471), .B(n2428), .O(n1065));
  andx g0967(.A(n1472), .B(pi00), .O(n1066));
  andx g0968(.A(n2647), .B(n2571), .O(n1067));
  andx g0969(.A(n1274), .B(pi05), .O(n1068));
  andx g0970(.A(n2378), .B(pi05), .O(n1069));
  andx g0971(.A(n2646), .B(n2573), .O(n1070));
  andx g0972(.A(n1474), .B(n2428), .O(n1071));
  andx g0973(.A(n1475), .B(pi00), .O(n1072));
  andx g0974(.A(n1473), .B(n2516), .O(n1073));
  andx g0975(.A(n1476), .B(pi04), .O(n1074));
  andx g0976(.A(n1479), .B(n1478), .O(n1075));
  andx g0977(.A(n1481), .B(n1480), .O(n1076));
  andx g0978(.A(n1483), .B(n1482), .O(n1077));
  andx g0979(.A(n1477), .B(n2362), .O(n1078));
  andx g0980(.A(n325), .B(pi06), .O(n1079));
  orx  g0981(.A(n169), .B(n2528), .O(n1080));
  orx  g0982(.A(n2368), .B(n2484), .O(n1081));
  orx  g0983(.A(n2459), .B(pi02), .O(n1082));
  orx  g0984(.A(n2671), .B(n168), .O(n1083));
  orx  g0985(.A(n171), .B(n170), .O(n1084));
  orx  g0986(.A(n173), .B(n2672), .O(n1085));
  orx  g0987(.A(n2672), .B(n2366), .O(n1086));
  orx  g0988(.A(n2585), .B(n174), .O(n1087));
  orx  g0989(.A(n283), .B(n2586), .O(n1088));
  orx  g0990(.A(n2383), .B(pi03), .O(n1089));
  orx  g0991(.A(n2626), .B(n2529), .O(n1090));
  orx  g0992(.A(n2626), .B(n2338), .O(n1091));
  orx  g0993(.A(n279), .B(n2528), .O(n1092));
  orx  g0994(.A(n2609), .B(n2585), .O(n1093));
  orx  g0995(.A(n2730), .B(n2586), .O(n1094));
  orx  g0996(.A(n177), .B(n2722), .O(n1095));
  orx  g0997(.A(n179), .B(n178), .O(n1096));
  orx  g0998(.A(n180), .B(n2626), .O(n1097));
  orx  g0999(.A(n333), .B(n334), .O(n1098));
  orx  g1000(.A(n337), .B(n338), .O(n1099));
  orx  g1001(.A(n339), .B(n340), .O(n1100));
  orx  g1002(.A(n343), .B(n344), .O(n1101));
  orx  g1003(.A(n345), .B(n346), .O(n1102));
  orx  g1004(.A(n347), .B(n348), .O(n1103));
  orx  g1005(.A(n349), .B(n350), .O(n1104));
  orx  g1006(.A(n2346), .B(n2440), .O(n1105));
  orx  g1007(.A(pi00), .B(n212), .O(n1106));
  orx  g1008(.A(n356), .B(n357), .O(n1107));
  orx  g1009(.A(n358), .B(n359), .O(n1108));
  orx  g1010(.A(n362), .B(n363), .O(n1109));
  orx  g1011(.A(n368), .B(n369), .O(n1110));
  orx  g1012(.A(n370), .B(n371), .O(n1111));
  orx  g1013(.A(n372), .B(n373), .O(n1112));
  orx  g1014(.A(n374), .B(n375), .O(n1113));
  orx  g1015(.A(n380), .B(n381), .O(n1114));
  orx  g1016(.A(n382), .B(n383), .O(n1115));
  orx  g1017(.A(n384), .B(n385), .O(n1116));
  orx  g1018(.A(pi04), .B(n2744), .O(n1117));
  orx  g1019(.A(n2500), .B(n388), .O(n1118));
  orx  g1020(.A(pi00), .B(n2663), .O(n1119));
  orx  g1021(.A(n2404), .B(n218), .O(n1120));
  orx  g1022(.A(pi04), .B(n392), .O(n1121));
  orx  g1023(.A(n2650), .B(n2528), .O(n1122));
  orx  g1024(.A(n400), .B(n401), .O(n1123));
  orx  g1025(.A(n406), .B(n407), .O(n1124));
  orx  g1026(.A(n408), .B(n409), .O(n1125));
  orx  g1027(.A(n412), .B(n413), .O(n1126));
  orx  g1028(.A(n414), .B(n415), .O(n1127));
  orx  g1029(.A(n416), .B(n417), .O(n1128));
  orx  g1030(.A(n2346), .B(n2442), .O(n1129));
  orx  g1031(.A(pi00), .B(n224), .O(n1130));
  orx  g1032(.A(n2663), .B(n2529), .O(n1131));
  orx  g1033(.A(pi04), .B(n420), .O(n1132));
  orx  g1034(.A(n428), .B(n429), .O(n1133));
  orx  g1035(.A(n434), .B(n435), .O(n1134));
  orx  g1036(.A(n436), .B(n437), .O(n1135));
  orx  g1037(.A(n438), .B(n439), .O(n1136));
  orx  g1038(.A(n442), .B(n443), .O(n1137));
  orx  g1039(.A(n444), .B(n445), .O(n1138));
  orx  g1040(.A(n446), .B(n447), .O(n1139));
  orx  g1041(.A(n448), .B(n449), .O(n1140));
  orx  g1042(.A(pi00), .B(n2662), .O(n1141));
  orx  g1043(.A(n2404), .B(n209), .O(n1142));
  orx  g1044(.A(n453), .B(n454), .O(n1143));
  orx  g1045(.A(n457), .B(n458), .O(n1144));
  orx  g1046(.A(n459), .B(n460), .O(n1145));
  orx  g1047(.A(n461), .B(n462), .O(n1146));
  orx  g1048(.A(n463), .B(n464), .O(n1147));
  orx  g1049(.A(n467), .B(n468), .O(n1148));
  orx  g1050(.A(n469), .B(n470), .O(n1149));
  orx  g1051(.A(n471), .B(n472), .O(n1150));
  orx  g1052(.A(pi04), .B(n2586), .O(n1151));
  orx  g1053(.A(n169), .B(n2528), .O(n1152));
  orx  g1054(.A(n2405), .B(n2608), .O(n1153));
  orx  g1055(.A(pi00), .B(n2640), .O(n1154));
  orx  g1056(.A(pi04), .B(n476), .O(n1155));
  orx  g1057(.A(n2607), .B(n2529), .O(n1156));
  orx  g1058(.A(n480), .B(n481), .O(n1157));
  orx  g1059(.A(n482), .B(n483), .O(n1158));
  orx  g1060(.A(n484), .B(n485), .O(n1159));
  orx  g1061(.A(n486), .B(n487), .O(n1160));
  orx  g1062(.A(n488), .B(n489), .O(n1161));
  orx  g1063(.A(n490), .B(n491), .O(n1162));
  orx  g1064(.A(n492), .B(n493), .O(n1163));
  orx  g1065(.A(n494), .B(n495), .O(n1164));
  orx  g1066(.A(n496), .B(n497), .O(n1165));
  orx  g1067(.A(pi00), .B(n2667), .O(n1166));
  orx  g1068(.A(n2729), .B(n2440), .O(n1167));
  orx  g1069(.A(pi00), .B(n244), .O(n1168));
  orx  g1070(.A(n2599), .B(n2765), .O(n1169));
  orx  g1071(.A(pi04), .B(n498), .O(n1170));
  orx  g1072(.A(n2501), .B(n501), .O(n1171));
  orx  g1073(.A(n505), .B(n506), .O(n1172));
  orx  g1074(.A(n507), .B(n508), .O(n1173));
  orx  g1075(.A(n509), .B(n510), .O(n1174));
  orx  g1076(.A(n511), .B(n512), .O(n1175));
  orx  g1077(.A(n513), .B(n514), .O(n1176));
  orx  g1078(.A(n517), .B(n518), .O(n1177));
  orx  g1079(.A(n519), .B(n520), .O(n1178));
  orx  g1080(.A(n521), .B(n522), .O(n1179));
  orx  g1081(.A(n523), .B(n524), .O(n1180));
  orx  g1082(.A(pi00), .B(n248), .O(n1181));
  orx  g1083(.A(n2665), .B(n2440), .O(n1182));
  orx  g1084(.A(n2405), .B(n2605), .O(n1183));
  orx  g1085(.A(pi00), .B(n2640), .O(n1184));
  orx  g1086(.A(pi04), .B(n527), .O(n1185));
  orx  g1087(.A(n2499), .B(n528), .O(n1186));
  orx  g1088(.A(n2331), .B(n2638), .O(n1187));
  orx  g1089(.A(pi06), .B(n2609), .O(n1188));
  orx  g1090(.A(n533), .B(n534), .O(n1189));
  orx  g1091(.A(n535), .B(n536), .O(n1190));
  orx  g1092(.A(n2541), .B(n2349), .O(n1191));
  orx  g1093(.A(pi05), .B(n537), .O(n1192));
  orx  g1094(.A(n2541), .B(n226), .O(n1193));
  orx  g1095(.A(pi05), .B(n237), .O(n1194));
  orx  g1096(.A(n2458), .B(n2370), .O(n1195));
  orx  g1097(.A(pi03), .B(n2392), .O(n1196));
  orx  g1098(.A(n541), .B(n542), .O(n1197));
  orx  g1099(.A(n543), .B(n544), .O(n1198));
  orx  g1100(.A(n545), .B(n546), .O(n1199));
  orx  g1101(.A(n549), .B(n550), .O(n1200));
  orx  g1102(.A(n551), .B(n552), .O(n1201));
  orx  g1103(.A(n554), .B(n555), .O(n1202));
  orx  g1104(.A(n556), .B(n557), .O(n1203));
  orx  g1105(.A(n558), .B(n559), .O(n1204));
  orx  g1106(.A(n560), .B(n561), .O(n1205));
  orx  g1107(.A(n562), .B(n563), .O(n1206));
  orx  g1108(.A(n564), .B(n565), .O(n1207));
  orx  g1109(.A(n566), .B(n567), .O(n1208));
  orx  g1110(.A(pi04), .B(n2674), .O(n1209));
  orx  g1111(.A(n2501), .B(n2643), .O(n1210));
  orx  g1112(.A(pi00), .B(n568), .O(n1211));
  orx  g1113(.A(n2405), .B(n257), .O(n1212));
  orx  g1114(.A(n574), .B(n575), .O(n1213));
  orx  g1115(.A(n576), .B(n577), .O(n1214));
  orx  g1116(.A(n578), .B(n579), .O(n1215));
  orx  g1117(.A(n580), .B(n581), .O(n1216));
  orx  g1118(.A(n585), .B(n586), .O(n1217));
  orx  g1119(.A(n589), .B(n590), .O(n1218));
  orx  g1120(.A(n591), .B(n592), .O(n1219));
  orx  g1121(.A(n593), .B(n594), .O(n1220));
  orx  g1122(.A(pi00), .B(n2398), .O(n1221));
  orx  g1123(.A(n2406), .B(n202), .O(n1222));
  orx  g1124(.A(n597), .B(n598), .O(n1223));
  orx  g1125(.A(n599), .B(n600), .O(n1224));
  orx  g1126(.A(n603), .B(n604), .O(n1225));
  orx  g1127(.A(n605), .B(n606), .O(n1226));
  orx  g1128(.A(n607), .B(n608), .O(n1227));
  orx  g1129(.A(n609), .B(n610), .O(n1228));
  orx  g1130(.A(n611), .B(n612), .O(n1229));
  orx  g1131(.A(n613), .B(n614), .O(n1230));
  orx  g1132(.A(n615), .B(n616), .O(n1231));
  orx  g1133(.A(n617), .B(n618), .O(n1232));
  orx  g1134(.A(n619), .B(n620), .O(n1233));
  orx  g1135(.A(n2404), .B(n2649), .O(n1234));
  orx  g1136(.A(pi00), .B(n244), .O(n1235));
  orx  g1137(.A(n2501), .B(n241), .O(n1236));
  orx  g1138(.A(pi04), .B(n621), .O(n1237));
  orx  g1139(.A(n625), .B(n626), .O(n1238));
  orx  g1140(.A(n627), .B(n628), .O(n1239));
  orx  g1141(.A(n629), .B(n630), .O(n1240));
  orx  g1142(.A(n631), .B(n632), .O(n1241));
  orx  g1143(.A(n633), .B(n634), .O(n1242));
  orx  g1144(.A(n637), .B(n638), .O(n1243));
  orx  g1145(.A(n639), .B(n640), .O(n1244));
  orx  g1146(.A(n641), .B(n642), .O(n1245));
  orx  g1147(.A(pi00), .B(n645), .O(n1246));
  orx  g1148(.A(n2406), .B(n267), .O(n1247));
  orx  g1149(.A(n651), .B(n652), .O(n1248));
  orx  g1150(.A(n653), .B(n654), .O(n1249));
  orx  g1151(.A(n657), .B(n658), .O(n1250));
  orx  g1152(.A(n659), .B(n660), .O(n1251));
  orx  g1153(.A(n663), .B(n664), .O(n1252));
  orx  g1154(.A(n665), .B(n666), .O(n1253));
  orx  g1155(.A(n667), .B(n668), .O(n1254));
  orx  g1156(.A(n669), .B(n670), .O(n1255));
  orx  g1157(.A(n671), .B(n672), .O(n1256));
  orx  g1158(.A(n673), .B(n674), .O(n1257));
  orx  g1159(.A(pi00), .B(n227), .O(n1258));
  orx  g1160(.A(n2406), .B(n236), .O(n1259));
  orx  g1161(.A(n677), .B(n678), .O(n1260));
  orx  g1162(.A(n679), .B(n680), .O(n1261));
  orx  g1163(.A(n684), .B(n685), .O(n1262));
  orx  g1164(.A(n690), .B(n691), .O(n1263));
  orx  g1165(.A(n692), .B(n693), .O(n1264));
  orx  g1166(.A(n694), .B(n695), .O(n1265));
  orx  g1167(.A(n696), .B(n697), .O(n1266));
  orx  g1168(.A(n698), .B(n699), .O(n1267));
  orx  g1169(.A(n700), .B(n701), .O(n1268));
  orx  g1170(.A(pi00), .B(n234), .O(n1269));
  orx  g1171(.A(n2407), .B(n274), .O(n1270));
  orx  g1172(.A(n705), .B(n706), .O(n1271));
  orx  g1173(.A(n707), .B(n708), .O(n1272));
  orx  g1174(.A(n712), .B(n713), .O(n1273));
  orx  g1175(.A(n714), .B(n715), .O(n1274));
  orx  g1176(.A(n716), .B(n717), .O(n1275));
  orx  g1177(.A(n718), .B(n719), .O(n1276));
  orx  g1178(.A(n720), .B(n721), .O(n1277));
  orx  g1179(.A(n722), .B(n723), .O(n1278));
  orx  g1180(.A(n724), .B(n725), .O(n1279));
  orx  g1181(.A(n726), .B(n727), .O(n1280));
  orx  g1182(.A(pi00), .B(n280), .O(n1281));
  orx  g1183(.A(n2405), .B(n279), .O(n1282));
  orx  g1184(.A(n733), .B(n734), .O(n1283));
  orx  g1185(.A(n735), .B(n736), .O(n1284));
  orx  g1186(.A(n739), .B(n740), .O(n1285));
  orx  g1187(.A(n741), .B(n742), .O(n1286));
  orx  g1188(.A(n743), .B(n744), .O(n1287));
  orx  g1189(.A(n747), .B(n748), .O(n1288));
  orx  g1190(.A(n751), .B(n752), .O(n1289));
  orx  g1191(.A(n753), .B(n754), .O(n1290));
  orx  g1192(.A(pi00), .B(n2727), .O(n1291));
  orx  g1193(.A(n2407), .B(n196), .O(n1292));
  orx  g1194(.A(pi00), .B(n2604), .O(n1293));
  orx  g1195(.A(n2662), .B(n2441), .O(n1294));
  orx  g1196(.A(pi04), .B(n755), .O(n1295));
  orx  g1197(.A(n2500), .B(n756), .O(n1296));
  orx  g1198(.A(n760), .B(n761), .O(n1297));
  orx  g1199(.A(n762), .B(n763), .O(n1298));
  orx  g1200(.A(n764), .B(n765), .O(n1299));
  orx  g1201(.A(n768), .B(n769), .O(n1300));
  orx  g1202(.A(n770), .B(n771), .O(n1301));
  orx  g1203(.A(n772), .B(n773), .O(n1302));
  orx  g1204(.A(n774), .B(n775), .O(n1303));
  orx  g1205(.A(n777), .B(n778), .O(n1304));
  orx  g1206(.A(n779), .B(n780), .O(n1305));
  orx  g1207(.A(n783), .B(n784), .O(n1306));
  orx  g1208(.A(n785), .B(n786), .O(n1307));
  orx  g1209(.A(n787), .B(n788), .O(n1308));
  orx  g1210(.A(n789), .B(n790), .O(n1309));
  orx  g1211(.A(n791), .B(n792), .O(n1310));
  orx  g1212(.A(n793), .B(n794), .O(n1311));
  orx  g1213(.A(n795), .B(n796), .O(n1312));
  orx  g1214(.A(n2459), .B(n2355), .O(n1313));
  orx  g1215(.A(pi02), .B(pi03), .O(n1314));
  orx  g1216(.A(pi00), .B(n199), .O(n1315));
  orx  g1217(.A(n2407), .B(n797), .O(n1316));
  orx  g1218(.A(n799), .B(n800), .O(n1317));
  orx  g1219(.A(n801), .B(n802), .O(n1318));
  orx  g1220(.A(n807), .B(n808), .O(n1319));
  orx  g1221(.A(n809), .B(n810), .O(n1320));
  orx  g1222(.A(n811), .B(n812), .O(n1321));
  orx  g1223(.A(n813), .B(n814), .O(n1322));
  orx  g1224(.A(n815), .B(n816), .O(n1323));
  orx  g1225(.A(n817), .B(n818), .O(n1324));
  orx  g1226(.A(n819), .B(n820), .O(n1325));
  orx  g1227(.A(n2458), .B(n2361), .O(n1326));
  orx  g1228(.A(pi03), .B(n2347), .O(n1327));
  orx  g1229(.A(n2406), .B(n189), .O(n1328));
  orx  g1230(.A(pi00), .B(n821), .O(n1329));
  orx  g1231(.A(n823), .B(n824), .O(n1330));
  orx  g1232(.A(n825), .B(n826), .O(n1331));
  orx  g1233(.A(n831), .B(n832), .O(n1332));
  orx  g1234(.A(n833), .B(n834), .O(n1333));
  orx  g1235(.A(n835), .B(n836), .O(n1334));
  orx  g1236(.A(n837), .B(n838), .O(n1335));
  orx  g1237(.A(n839), .B(n840), .O(n1336));
  orx  g1238(.A(n841), .B(n842), .O(n1337));
  orx  g1239(.A(pi04), .B(n187), .O(n1338));
  orx  g1240(.A(n2500), .B(n228), .O(n1339));
  orx  g1241(.A(pi00), .B(n843), .O(n1340));
  orx  g1242(.A(n2408), .B(n844), .O(n1341));
  orx  g1243(.A(n848), .B(n849), .O(n1342));
  orx  g1244(.A(n850), .B(n851), .O(n1343));
  orx  g1245(.A(n852), .B(n853), .O(n1344));
  orx  g1246(.A(n854), .B(n855), .O(n1345));
  orx  g1247(.A(n857), .B(n858), .O(n1346));
  orx  g1248(.A(n859), .B(n860), .O(n1347));
  orx  g1249(.A(n861), .B(n862), .O(n1348));
  orx  g1250(.A(pi00), .B(n167), .O(n1349));
  orx  g1251(.A(n2408), .B(n299), .O(n1350));
  orx  g1252(.A(n2408), .B(n2643), .O(n1351));
  orx  g1253(.A(pi00), .B(n2640), .O(n1352));
  orx  g1254(.A(pi04), .B(n865), .O(n1353));
  orx  g1255(.A(n2502), .B(n866), .O(n1354));
  orx  g1256(.A(n870), .B(n871), .O(n1355));
  orx  g1257(.A(n872), .B(n873), .O(n1356));
  orx  g1258(.A(n874), .B(n875), .O(n1357));
  orx  g1259(.A(n876), .B(n877), .O(n1358));
  orx  g1260(.A(n878), .B(n879), .O(n1359));
  orx  g1261(.A(n880), .B(n881), .O(n1360));
  orx  g1262(.A(pi04), .B(n229), .O(n1361));
  orx  g1263(.A(n2496), .B(n2640), .O(n1362));
  orx  g1264(.A(pi00), .B(n882), .O(n1363));
  orx  g1265(.A(n2407), .B(n302), .O(n1364));
  orx  g1266(.A(n886), .B(n887), .O(n1365));
  orx  g1267(.A(n888), .B(n889), .O(n1366));
  orx  g1268(.A(n890), .B(n891), .O(n1367));
  orx  g1269(.A(n892), .B(n893), .O(n1368));
  orx  g1270(.A(n894), .B(n895), .O(n1369));
  orx  g1271(.A(n2409), .B(n2637), .O(n1370));
  orx  g1272(.A(pi00), .B(n200), .O(n1371));
  orx  g1273(.A(n897), .B(n898), .O(n1372));
  orx  g1274(.A(n899), .B(n900), .O(n1373));
  orx  g1275(.A(n903), .B(n904), .O(n1374));
  orx  g1276(.A(n905), .B(n906), .O(n1375));
  orx  g1277(.A(n907), .B(n908), .O(n1376));
  orx  g1278(.A(n909), .B(n910), .O(n1377));
  orx  g1279(.A(n911), .B(n912), .O(n1378));
  orx  g1280(.A(n913), .B(n914), .O(n1379));
  orx  g1281(.A(n915), .B(n916), .O(n1380));
  orx  g1282(.A(n917), .B(n918), .O(n1381));
  orx  g1283(.A(n919), .B(n920), .O(n1382));
  orx  g1284(.A(n923), .B(n924), .O(n1383));
  orx  g1285(.A(n925), .B(n926), .O(n1384));
  orx  g1286(.A(n927), .B(n928), .O(n1385));
  orx  g1287(.A(n929), .B(n930), .O(n1386));
  orx  g1288(.A(n931), .B(n932), .O(n1387));
  orx  g1289(.A(n933), .B(n934), .O(n1388));
  orx  g1290(.A(n935), .B(n936), .O(n1389));
  orx  g1291(.A(n2409), .B(n553), .O(n1390));
  orx  g1292(.A(pi00), .B(n2616), .O(n1391));
  orx  g1293(.A(n938), .B(n939), .O(n1392));
  orx  g1294(.A(n942), .B(n943), .O(n1393));
  orx  g1295(.A(n944), .B(n945), .O(n1394));
  orx  g1296(.A(n946), .B(n947), .O(n1395));
  orx  g1297(.A(n948), .B(n949), .O(n1396));
  orx  g1298(.A(n950), .B(n951), .O(n1397));
  orx  g1299(.A(n952), .B(n953), .O(n1398));
  orx  g1300(.A(n954), .B(n955), .O(n1399));
  orx  g1301(.A(n956), .B(n957), .O(n1400));
  orx  g1302(.A(pi00), .B(n2528), .O(n1401));
  orx  g1303(.A(pi04), .B(n2586), .O(n1402));
  orx  g1304(.A(pi00), .B(n200), .O(n1403));
  orx  g1305(.A(n2409), .B(n211), .O(n1404));
  orx  g1306(.A(n2617), .B(n2529), .O(n1405));
  orx  g1307(.A(pi04), .B(n959), .O(n1406));
  orx  g1308(.A(n965), .B(n966), .O(n1407));
  orx  g1309(.A(n967), .B(n968), .O(n1408));
  orx  g1310(.A(n969), .B(n970), .O(n1409));
  orx  g1311(.A(n971), .B(n972), .O(n1410));
  orx  g1312(.A(n973), .B(n974), .O(n1411));
  orx  g1313(.A(n975), .B(n976), .O(n1412));
  orx  g1314(.A(n977), .B(n978), .O(n1413));
  orx  g1315(.A(n979), .B(n980), .O(n1414));
  orx  g1316(.A(pi00), .B(n2645), .O(n1415));
  orx  g1317(.A(n2403), .B(n267), .O(n1416));
  orx  g1318(.A(n982), .B(n983), .O(n1417));
  orx  g1319(.A(n986), .B(n987), .O(n1418));
  orx  g1320(.A(n988), .B(n989), .O(n1419));
  orx  g1321(.A(n990), .B(n991), .O(n1420));
  orx  g1322(.A(n992), .B(n993), .O(n1421));
  orx  g1323(.A(n994), .B(n995), .O(n1422));
  orx  g1324(.A(n996), .B(n997), .O(n1423));
  orx  g1325(.A(pi03), .B(n2387), .O(n1424));
  orx  g1326(.A(n2458), .B(n2368), .O(n1425));
  orx  g1327(.A(pi00), .B(n2671), .O(n1426));
  orx  g1328(.A(n2409), .B(n998), .O(n1427));
  orx  g1329(.A(n2730), .B(n2440), .O(n1428));
  orx  g1330(.A(pi00), .B(n279), .O(n1429));
  orx  g1331(.A(pi04), .B(n999), .O(n1430));
  orx  g1332(.A(n2502), .B(n1000), .O(n1431));
  orx  g1333(.A(n1004), .B(n1005), .O(n1432));
  orx  g1334(.A(n1006), .B(n1007), .O(n1433));
  orx  g1335(.A(n1008), .B(n1009), .O(n1434));
  orx  g1336(.A(n1010), .B(n1011), .O(n1435));
  orx  g1337(.A(n1012), .B(n1013), .O(n1436));
  orx  g1338(.A(n1014), .B(n1015), .O(n1437));
  orx  g1339(.A(n1016), .B(n1017), .O(n1438));
  orx  g1340(.A(n2729), .B(n2442), .O(n1439));
  orx  g1341(.A(pi00), .B(n2618), .O(n1440));
  orx  g1342(.A(pi00), .B(n2643), .O(n1441));
  orx  g1343(.A(n2408), .B(n248), .O(n1442));
  orx  g1344(.A(pi04), .B(n1018), .O(n1443));
  orx  g1345(.A(n2502), .B(n1019), .O(n1444));
  orx  g1346(.A(n1023), .B(n1024), .O(n1445));
  orx  g1347(.A(n1025), .B(n1026), .O(n1446));
  orx  g1348(.A(n1027), .B(n1028), .O(n1447));
  orx  g1349(.A(n1029), .B(n1030), .O(n1448));
  orx  g1350(.A(n1031), .B(n1032), .O(n1449));
  orx  g1351(.A(n1033), .B(n1034), .O(n1450));
  orx  g1352(.A(n1035), .B(n1036), .O(n1451));
  orx  g1353(.A(n1037), .B(n1038), .O(n1452));
  orx  g1354(.A(n2500), .B(n244), .O(n1453));
  orx  g1355(.A(pi04), .B(n315), .O(n1454));
  orx  g1356(.A(pi04), .B(n240), .O(n1455));
  orx  g1357(.A(n2597), .B(n2529), .O(n1456));
  orx  g1358(.A(pi00), .B(n1039), .O(n1457));
  orx  g1359(.A(n2410), .B(n1040), .O(n1458));
  orx  g1360(.A(n1044), .B(n1045), .O(n1459));
  orx  g1361(.A(n1046), .B(n1047), .O(n1460));
  orx  g1362(.A(n1048), .B(n1049), .O(n1461));
  orx  g1363(.A(n1050), .B(n1051), .O(n1462));
  orx  g1364(.A(n1052), .B(n1053), .O(n1463));
  orx  g1365(.A(n1054), .B(n1055), .O(n1464));
  orx  g1366(.A(pi04), .B(n2633), .O(n1465));
  orx  g1367(.A(n2502), .B(n2612), .O(n1466));
  orx  g1368(.A(n2730), .B(n2527), .O(n1467));
  orx  g1369(.A(pi04), .B(n2668), .O(n1468));
  orx  g1370(.A(pi00), .B(n1056), .O(n1469));
  orx  g1371(.A(n2410), .B(n1057), .O(n1470));
  orx  g1372(.A(n1061), .B(n1062), .O(n1471));
  orx  g1373(.A(n1063), .B(n1064), .O(n1472));
  orx  g1374(.A(n1065), .B(n1066), .O(n1473));
  orx  g1375(.A(n1067), .B(n1068), .O(n1474));
  orx  g1376(.A(n1069), .B(n1070), .O(n1475));
  orx  g1377(.A(n1071), .B(n1072), .O(n1476));
  orx  g1378(.A(n1073), .B(n1074), .O(n1477));
  orx  g1379(.A(n2602), .B(n2441), .O(n1478));
  orx  g1380(.A(pi00), .B(n2613), .O(n1479));
  orx  g1381(.A(pi00), .B(n2603), .O(n1480));
  orx  g1382(.A(n2663), .B(n2441), .O(n1481));
  orx  g1383(.A(pi04), .B(n1075), .O(n1482));
  orx  g1384(.A(n2501), .B(n1076), .O(n1483));
  orx  g1385(.A(n2330), .B(pi01), .O(n1484));
  orx  g1386(.A(pi02), .B(pi01), .O(n1485));
  orx  g1387(.A(n2390), .B(n2701), .O(n1486));
  orx  g1388(.A(n2389), .B(pi00), .O(n1487));
  andx g1389(.A(n2150), .B(pi05), .O(n1488));
  orx  g1390(.A(n2379), .B(n2441), .O(n1489));
  andx g1391(.A(n1489), .B(pi04), .O(n1490));
  orx  g1392(.A(n1504), .B(n2442), .O(n1491));
  andx g1393(.A(n2698), .B(pi04), .O(n1492));
  andx g1394(.A(n2366), .B(n2430), .O(n1493));
  orx  g1395(.A(n2710), .B(n2382), .O(n1494));
  andx g1396(.A(pi05), .B(n2726), .O(n1495));
  orx  g1397(.A(n2388), .B(n2485), .O(n1496));
  orx  g1398(.A(n1505), .B(pi03), .O(n1497));
  andx g1399(.A(n2037), .B(n2677), .O(n1498));
  orx  g1400(.A(pi05), .B(pi04), .O(n1499));
  orx  g1401(.A(n2706), .B(n2366), .O(n1500));
  orx  g1402(.A(n2719), .B(n2371), .O(n1501));
  orx  g1403(.A(n2718), .B(n2689), .O(n1502));
  orx  g1404(.A(n2340), .B(n2689), .O(n1503));
  orx  g1405(.A(n2361), .B(n2356), .O(n1504));
  orx  g1406(.A(pi00), .B(n2380), .O(n1505));
  orx  g1407(.A(n2498), .B(n2485), .O(n1506));
  orx  g1408(.A(pi00), .B(n2371), .O(n1507));
  andx g1409(.A(n1591), .B(n2471), .O(n1508));
  andx g1410(.A(n2585), .B(n2048), .O(n1509));
  andx g1411(.A(n2681), .B(n1555), .O(n1510));
  orx  g1412(.A(n1600), .B(n1601), .O(n1511));
  orx  g1413(.A(n1669), .B(n1670), .O(n1512));
  orx  g1414(.A(n1655), .B(n1656), .O(n1513));
  orx  g1415(.A(n1732), .B(n1733), .O(n1514));
  orx  g1416(.A(n1906), .B(n1907), .O(n1515));
  orx  g1417(.A(n1888), .B(n1887), .O(n1516));
  orx  g1418(.A(n1948), .B(n1949), .O(n1517));
  orx  g1419(.A(n2007), .B(n2008), .O(n1518));
  orx  g1420(.A(n1614), .B(n1615), .O(n1519));
  andx g1421(.A(n1617), .B(n2516), .O(n1520));
  andx g1422(.A(n1618), .B(n2574), .O(n1521));
  orx  g1423(.A(n1620), .B(n1619), .O(n1522));
  orx  g1424(.A(n1635), .B(n1636), .O(n1523));
  orx  g1425(.A(n1625), .B(n1626), .O(n1524));
  andx g1426(.A(n1646), .B(n2574), .O(n1525));
  orx  g1427(.A(n1648), .B(n1647), .O(n1526));
  andx g1428(.A(n2394), .B(n2517), .O(n1527));
  andx g1429(.A(n1672), .B(n2572), .O(n1528));
  orx  g1430(.A(n1674), .B(n1673), .O(n1529));
  orx  g1431(.A(n1698), .B(n1699), .O(n1530));
  andx g1432(.A(n1590), .B(n1702), .O(n1531));
  orx  g1433(.A(n1704), .B(n1703), .O(n1532));
  orx  g1434(.A(n1725), .B(n1726), .O(n1533));
  andx g1435(.A(n1519), .B(n2336), .O(n1534));
  orx  g1436(.A(n1711), .B(n1712), .O(n1535));
  andx g1437(.A(n1727), .B(n2351), .O(n1536));
  orx  g1438(.A(n1728), .B(n1729), .O(n1537));
  andx g1439(.A(n1750), .B(n1748), .O(n1538));
  orx  g1440(.A(n1752), .B(n1751), .O(n1539));
  orx  g1441(.A(n1761), .B(n1762), .O(n1540));
  orx  g1442(.A(n1755), .B(n1756), .O(n1541));
  andx g1443(.A(n1774), .B(n2574), .O(n1542));
  orx  g1444(.A(n1776), .B(n1775), .O(n1543));
  andx g1445(.A(n2380), .B(n2048), .O(n1544));
  andx g1446(.A(n1789), .B(n2062), .O(n1545));
  andx g1447(.A(n2061), .B(n2049), .O(n1546));
  orx  g1448(.A(n1777), .B(n1778), .O(n1547));
  andx g1449(.A(n1791), .B(n2575), .O(n1548));
  orx  g1450(.A(n1793), .B(n1792), .O(n1549));
  orx  g1451(.A(n1812), .B(n1813), .O(n1550));
  andx g1452(.A(n2365), .B(n1588), .O(n1551));
  andx g1453(.A(n1816), .B(n2573), .O(n1552));
  orx  g1454(.A(n1818), .B(n1817), .O(n1553));
  orx  g1455(.A(n1834), .B(n1835), .O(n1554));
  orx  g1456(.A(n1822), .B(n1823), .O(n1555));
  andx g1457(.A(n2063), .B(n1505), .O(n1556));
  andx g1458(.A(n1839), .B(n2575), .O(n1557));
  orx  g1459(.A(n1841), .B(n1840), .O(n1558));
  andx g1460(.A(n1864), .B(n2572), .O(n1559));
  orx  g1461(.A(n1866), .B(n1865), .O(n1560));
  andx g1462(.A(n1882), .B(n2573), .O(n1561));
  orx  g1463(.A(n1884), .B(n1883), .O(n1562));
  orx  g1464(.A(n1903), .B(n1904), .O(n1563));
  andx g1465(.A(n1909), .B(n2362), .O(n1564));
  orx  g1466(.A(n1910), .B(n1911), .O(n1565));
  orx  g1467(.A(n1912), .B(n1913), .O(n1566));
  andx g1468(.A(n1932), .B(n1929), .O(n1567));
  orx  g1469(.A(n1934), .B(n1933), .O(n1568));
  andx g1470(.A(n1951), .B(n2349), .O(n1569));
  orx  g1471(.A(n1952), .B(n1953), .O(n1570));
  andx g1472(.A(n2067), .B(n1491), .O(n1571));
  andx g1473(.A(n1971), .B(n2576), .O(n1572));
  orx  g1474(.A(n1973), .B(n1972), .O(n1573));
  andx g1475(.A(n1990), .B(n2576), .O(n1574));
  orx  g1476(.A(n1992), .B(n1991), .O(n1575));
  orx  g1477(.A(n2009), .B(n2010), .O(n1576));
  andx g1478(.A(n2068), .B(n2573), .O(n1577));
  orx  g1479(.A(n2012), .B(n2011), .O(n1578));
  andx g1480(.A(pi00), .B(pi02), .O(n1579));
  andx g1481(.A(n2070), .B(n2577), .O(n1580));
  orx  g1482(.A(n2026), .B(n2025), .O(n1581));
  andx g1483(.A(pi04), .B(n1497), .O(n1582));
  andx g1484(.A(n2071), .B(n2577), .O(n1583));
  orx  g1485(.A(n2036), .B(n2035), .O(n1584));
  orx  g1486(.A(n2040), .B(n2039), .O(n1585));
  orx  g1487(.A(n2041), .B(n2042), .O(n1586));
  orx  g1488(.A(n2043), .B(n2044), .O(n1587));
  orx  g1489(.A(n2332), .B(n2442), .O(n1588));
  orx  g1490(.A(n2718), .B(n2696), .O(n1589));
  andx g1491(.A(n1506), .B(n2574), .O(n1590));
  andx g1492(.A(n2585), .B(n2361), .O(n1591));
  andx g1493(.A(pi00), .B(n2359), .O(n1592));
  andx g1494(.A(n2718), .B(n2436), .O(n1593));
  andx g1495(.A(pi01), .B(n2430), .O(n1594));
  andx g1496(.A(pi00), .B(n2394), .O(n1595));
  andx g1497(.A(n2075), .B(n2517), .O(n1596));
  andx g1498(.A(n2076), .B(pi04), .O(n1597));
  andx g1499(.A(pi02), .B(n2434), .O(n1598));
  andx g1500(.A(pi00), .B(n2395), .O(n1599));
  andx g1501(.A(pi01), .B(n2358), .O(n1600));
  andx g1502(.A(pi02), .B(n2356), .O(n1601));
  andx g1503(.A(n2078), .B(n2518), .O(n1602));
  andx g1504(.A(n2726), .B(pi04), .O(n1603));
  andx g1505(.A(n2077), .B(n2472), .O(n1604));
  andx g1506(.A(n2079), .B(pi03), .O(n1605));
  andx g1507(.A(n2723), .B(n2518), .O(n1606));
  andx g1508(.A(n2724), .B(pi04), .O(n1607));
  andx g1509(.A(n1486), .B(n2517), .O(n1608));
  andx g1510(.A(n2725), .B(pi04), .O(n1609));
  andx g1511(.A(n2081), .B(n2471), .O(n1610));
  andx g1512(.A(n2082), .B(pi03), .O(n1611));
  andx g1513(.A(n2080), .B(n2578), .O(n1612));
  andx g1514(.A(n2083), .B(pi05), .O(n1613));
  andx g1515(.A(pi00), .B(pi02), .O(n1614));
  andx g1516(.A(n2365), .B(n2430), .O(n1615));
  andx g1517(.A(n2086), .B(n2085), .O(n1616));
  andx g1518(.A(n2088), .B(n2087), .O(n1617));
  andx g1519(.A(n2090), .B(n2089), .O(n1618));
  andx g1520(.A(n2084), .B(n2362), .O(n1619));
  andx g1521(.A(n1521), .B(pi06), .O(n1620));
  andx g1522(.A(pi04), .B(n2330), .O(n1621));
  andx g1523(.A(n2052), .B(n2519), .O(n1622));
  andx g1524(.A(pi00), .B(n2354), .O(n1623));
  andx g1525(.A(pi01), .B(n2431), .O(n1624));
  andx g1526(.A(pi02), .B(n2429), .O(n1625));
  andx g1527(.A(n2381), .B(pi00), .O(n1626));
  andx g1528(.A(n2092), .B(n2518), .O(n1627));
  andx g1529(.A(n1524), .B(pi04), .O(n1628));
  andx g1530(.A(n2091), .B(n2472), .O(n1629));
  andx g1531(.A(n2093), .B(pi03), .O(n1630));
  andx g1532(.A(pi02), .B(n2431), .O(n1631));
  andx g1533(.A(pi00), .B(n2390), .O(n1632));
  andx g1534(.A(n2051), .B(pi04), .O(n1633));
  andx g1535(.A(n2095), .B(n2520), .O(n1634));
  andx g1536(.A(pi02), .B(n2435), .O(n1635));
  andx g1537(.A(pi00), .B(n2344), .O(n1636));
  andx g1538(.A(n1487), .B(n2519), .O(n1637));
  andx g1539(.A(n1523), .B(pi04), .O(n1638));
  andx g1540(.A(n2096), .B(n2472), .O(n1639));
  andx g1541(.A(n2097), .B(pi03), .O(n1640));
  andx g1542(.A(n2094), .B(n2575), .O(n1641));
  andx g1543(.A(n2098), .B(pi05), .O(n1642));
  orx  g1544(.A(n2718), .B(n2441), .O(n1643));
  andx g1545(.A(n2101), .B(n2100), .O(n1644));
  andx g1546(.A(n2103), .B(n2102), .O(n1645));
  andx g1547(.A(n2105), .B(n2104), .O(n1646));
  andx g1548(.A(n2099), .B(n2353), .O(n1647));
  andx g1549(.A(n1525), .B(pi06), .O(n1648));
  andx g1550(.A(pi01), .B(n2427), .O(n1649));
  andx g1551(.A(n2333), .B(pi00), .O(n1650));
  andx g1552(.A(n1502), .B(n2520), .O(n1651));
  andx g1553(.A(n2106), .B(pi04), .O(n1652));
  andx g1554(.A(n2390), .B(n2525), .O(n1653));
  andx g1555(.A(pi04), .B(n1504), .O(n1654));
  andx g1556(.A(pi00), .B(n2519), .O(n1655));
  andx g1557(.A(pi04), .B(n2432), .O(n1656));
  andx g1558(.A(n1513), .B(pi01), .O(n1657));
  andx g1559(.A(n2108), .B(n2679), .O(n1658));
  andx g1560(.A(n2107), .B(n2473), .O(n1659));
  andx g1561(.A(n2109), .B(pi03), .O(n1660));
  andx g1562(.A(n2395), .B(n2429), .O(n1661));
  andx g1563(.A(n2373), .B(pi00), .O(n1662));
  andx g1564(.A(n2053), .B(n2505), .O(n1663));
  andx g1565(.A(n2111), .B(pi04), .O(n1664));
  andx g1566(.A(n2112), .B(n2472), .O(n1665));
  andx g1567(.A(n2054), .B(pi03), .O(n1666));
  andx g1568(.A(n2110), .B(n2578), .O(n1667));
  andx g1569(.A(n2113), .B(pi05), .O(n1668));
  andx g1570(.A(n2332), .B(pi00), .O(n1669));
  andx g1571(.A(n2382), .B(n2432), .O(n1670));
  andx g1572(.A(n2116), .B(n2115), .O(n1671));
  andx g1573(.A(n2118), .B(n2117), .O(n1672));
  andx g1574(.A(n2114), .B(n2335), .O(n1673));
  andx g1575(.A(n1528), .B(pi06), .O(n1674));
  andx g1576(.A(n2382), .B(n2431), .O(n1675));
  andx g1577(.A(pi00), .B(n2389), .O(n1676));
  andx g1578(.A(pi00), .B(n2359), .O(n1677));
  andx g1579(.A(n2393), .B(n2429), .O(n1678));
  andx g1580(.A(n2119), .B(n2578), .O(n1679));
  andx g1581(.A(n2120), .B(pi05), .O(n1680));
  andx g1582(.A(pi05), .B(pi00), .O(n1681));
  andx g1583(.A(n2055), .B(n2576), .O(n1682));
  andx g1584(.A(n2121), .B(n2473), .O(n1683));
  andx g1585(.A(n2122), .B(pi03), .O(n1684));
  andx g1586(.A(pi00), .B(pi02), .O(n1685));
  andx g1587(.A(n2385), .B(n2433), .O(n1686));
  andx g1588(.A(n2056), .B(n2579), .O(n1687));
  andx g1589(.A(n2124), .B(pi05), .O(n1688));
  andx g1590(.A(n2333), .B(n2430), .O(n1689));
  andx g1591(.A(pi00), .B(n2343), .O(n1690));
  andx g1592(.A(n2128), .B(n2127), .O(n1691));
  andx g1593(.A(n2126), .B(n2579), .O(n1692));
  andx g1594(.A(n1691), .B(pi05), .O(n1693));
  andx g1595(.A(n2125), .B(n2473), .O(n1694));
  andx g1596(.A(n2129), .B(pi03), .O(n1695));
  andx g1597(.A(n2123), .B(n2520), .O(n1696));
  andx g1598(.A(n2130), .B(pi04), .O(n1697));
  andx g1599(.A(n2355), .B(n2434), .O(n1698));
  andx g1600(.A(pi00), .B(n2388), .O(n1699));
  orx  g1601(.A(pi00), .B(n2365), .O(n1700));
  andx g1602(.A(n2133), .B(n2132), .O(n1701));
  andx g1603(.A(n2135), .B(n2134), .O(n1702));
  andx g1604(.A(n2131), .B(n2336), .O(n1703));
  andx g1605(.A(n1531), .B(pi06), .O(n1704));
  andx g1606(.A(pi02), .B(n2432), .O(n1705));
  andx g1607(.A(n2332), .B(pi00), .O(n1706));
  andx g1608(.A(n2124), .B(n2363), .O(n1707));
  andx g1609(.A(n2136), .B(pi06), .O(n1708));
  andx g1610(.A(pi00), .B(pi02), .O(n1709));
  andx g1611(.A(n2381), .B(n2434), .O(n1710));
  andx g1612(.A(pi00), .B(pi01), .O(n1711));
  andx g1613(.A(n2340), .B(n2433), .O(n1712));
  andx g1614(.A(n2138), .B(n2352), .O(n1713));
  andx g1615(.A(n1535), .B(pi06), .O(n1714));
  andx g1616(.A(n2137), .B(n2474), .O(n1715));
  andx g1617(.A(n2139), .B(pi03), .O(n1716));
  andx g1618(.A(pi06), .B(n1500), .O(n1717));
  andx g1619(.A(n2719), .B(n2331), .O(n1718));
  andx g1620(.A(n2141), .B(n2474), .O(n1719));
  andx g1621(.A(n1534), .B(pi03), .O(n1720));
  andx g1622(.A(n2140), .B(n2503), .O(n1721));
  andx g1623(.A(n2142), .B(pi04), .O(n1722));
  andx g1624(.A(n2145), .B(n2144), .O(n1723));
  andx g1625(.A(n2147), .B(n2146), .O(n1724));
  andx g1626(.A(pi03), .B(pi04), .O(n1725));
  andx g1627(.A(pi00), .B(n2518), .O(n1726));
  andx g1628(.A(n2149), .B(n2148), .O(n1727));
  andx g1629(.A(n2143), .B(n2575), .O(n1728));
  andx g1630(.A(n1536), .B(pi05), .O(n1729));
  andx g1631(.A(pi00), .B(n2393), .O(n1730));
  andx g1632(.A(n2379), .B(n2435), .O(n1731));
  andx g1633(.A(n2380), .B(pi00), .O(n1732));
  andx g1634(.A(n2389), .B(n2431), .O(n1733));
  andx g1635(.A(n2356), .B(n2429), .O(n1734));
  andx g1636(.A(pi00), .B(n2394), .O(n1735));
  andx g1637(.A(n1514), .B(n2580), .O(n1736));
  andx g1638(.A(n2151), .B(pi05), .O(n1737));
  andx g1639(.A(n2057), .B(n2474), .O(n1738));
  andx g1640(.A(n2152), .B(pi03), .O(n1739));
  andx g1641(.A(pi05), .B(n2380), .O(n1740));
  andx g1642(.A(n1512), .B(n2580), .O(n1741));
  andx g1643(.A(pi05), .B(n2045), .O(n1742));
  andx g1644(.A(n2058), .B(n2577), .O(n1743));
  andx g1645(.A(n2154), .B(n2474), .O(n1744));
  andx g1646(.A(n2155), .B(pi03), .O(n1745));
  andx g1647(.A(n2153), .B(n2527), .O(n1746));
  andx g1648(.A(n2156), .B(pi04), .O(n1747));
  andx g1649(.A(n2159), .B(n2158), .O(n1748));
  andx g1650(.A(n2161), .B(n2160), .O(n1749));
  andx g1651(.A(n2163), .B(n2162), .O(n1750));
  andx g1652(.A(n2157), .B(n2336), .O(n1751));
  andx g1653(.A(n1538), .B(pi06), .O(n1752));
  andx g1654(.A(n2693), .B(pi04), .O(n1753));
  andx g1655(.A(n2690), .B(n2526), .O(n1754));
  andx g1656(.A(pi00), .B(pi01), .O(n1755));
  andx g1657(.A(n2372), .B(n2434), .O(n1756));
  andx g1658(.A(pi04), .B(n2436), .O(n1757));
  andx g1659(.A(n1541), .B(n2517), .O(n1758));
  andx g1660(.A(n2164), .B(n2475), .O(n1759));
  andx g1661(.A(n2165), .B(pi03), .O(n1760));
  andx g1662(.A(pi01), .B(n2434), .O(n1761));
  andx g1663(.A(n2342), .B(pi00), .O(n1762));
  andx g1664(.A(pi00), .B(n2358), .O(n1763));
  andx g1665(.A(n2341), .B(n2436), .O(n1764));
  andx g1666(.A(n2714), .B(pi04), .O(n1765));
  andx g1667(.A(n2167), .B(n2524), .O(n1766));
  andx g1668(.A(n2059), .B(n2475), .O(n1767));
  andx g1669(.A(n2168), .B(pi03), .O(n1768));
  andx g1670(.A(n2166), .B(n2580), .O(n1769));
  andx g1671(.A(n2169), .B(pi05), .O(n1770));
  orx  g1672(.A(n2689), .B(n2383), .O(n1771));
  andx g1673(.A(n2172), .B(n2171), .O(n1772));
  andx g1674(.A(n2174), .B(n2173), .O(n1773));
  andx g1675(.A(n2176), .B(n2175), .O(n1774));
  andx g1676(.A(n2170), .B(n2335), .O(n1775));
  andx g1677(.A(n1542), .B(pi06), .O(n1776));
  andx g1678(.A(pi00), .B(pi02), .O(n1777));
  andx g1679(.A(n2379), .B(n2433), .O(n1778));
  andx g1680(.A(n1502), .B(n2521), .O(n1779));
  andx g1681(.A(n1547), .B(pi04), .O(n1780));
  andx g1682(.A(n2177), .B(n2475), .O(n1781));
  andx g1683(.A(n2060), .B(pi03), .O(n1782));
  andx g1684(.A(pi04), .B(n2390), .O(n1783));
  andx g1685(.A(n2692), .B(n2519), .O(n1784));
  andx g1686(.A(n2179), .B(n2476), .O(n1785));
  andx g1687(.A(n1546), .B(pi03), .O(n1786));
  andx g1688(.A(n2178), .B(n2581), .O(n1787));
  andx g1689(.A(n2180), .B(pi05), .O(n1788));
  andx g1690(.A(n2183), .B(n2182), .O(n1789));
  andx g1691(.A(n2185), .B(n2184), .O(n1790));
  andx g1692(.A(n2187), .B(n2186), .O(n1791));
  andx g1693(.A(n2181), .B(n2351), .O(n1792));
  andx g1694(.A(n1548), .B(pi06), .O(n1793));
  andx g1695(.A(n2052), .B(n2578), .O(n1794));
  andx g1696(.A(n1551), .B(pi05), .O(n1795));
  andx g1697(.A(pi00), .B(n2718), .O(n1796));
  andx g1698(.A(n2340), .B(n2437), .O(n1797));
  andx g1699(.A(n2708), .B(pi05), .O(n1798));
  andx g1700(.A(n2189), .B(n2581), .O(n1799));
  andx g1701(.A(n2188), .B(n2475), .O(n1800));
  andx g1702(.A(n2190), .B(pi03), .O(n1801));
  andx g1703(.A(pi05), .B(n2435), .O(n1802));
  andx g1704(.A(pi02), .B(n2577), .O(n1803));
  andx g1705(.A(pi00), .B(pi01), .O(n1804));
  andx g1706(.A(n2394), .B(n2437), .O(n1805));
  andx g1707(.A(n1519), .B(n2579), .O(n1806));
  andx g1708(.A(n2193), .B(pi05), .O(n1807));
  andx g1709(.A(n2192), .B(n2476), .O(n1808));
  andx g1710(.A(n2194), .B(pi03), .O(n1809));
  andx g1711(.A(n2191), .B(n2522), .O(n1810));
  andx g1712(.A(n2195), .B(pi04), .O(n1811));
  andx g1713(.A(n2388), .B(n2435), .O(n1812));
  andx g1714(.A(n2342), .B(pi00), .O(n1813));
  andx g1715(.A(n2198), .B(n2197), .O(n1814));
  andx g1716(.A(n2200), .B(n2199), .O(n1815));
  andx g1717(.A(n2202), .B(n2201), .O(n1816));
  andx g1718(.A(n2196), .B(n2363), .O(n1817));
  andx g1719(.A(n1552), .B(pi06), .O(n1818));
  andx g1720(.A(n1489), .B(pi04), .O(n1819));
  andx g1721(.A(n1556), .B(n2477), .O(n1820));
  andx g1722(.A(n2203), .B(pi03), .O(n1821));
  andx g1723(.A(pi02), .B(n2438), .O(n1822));
  andx g1724(.A(n2380), .B(pi00), .O(n1823));
  andx g1725(.A(pi00), .B(n2392), .O(n1824));
  andx g1726(.A(n2718), .B(n2433), .O(n1825));
  andx g1727(.A(n2333), .B(pi00), .O(n1826));
  andx g1728(.A(n2343), .B(n2438), .O(n1827));
  andx g1729(.A(n2205), .B(n2522), .O(n1828));
  andx g1730(.A(n2206), .B(pi04), .O(n1829));
  andx g1731(.A(n2064), .B(n2477), .O(n1830));
  andx g1732(.A(n2207), .B(pi03), .O(n1831));
  andx g1733(.A(n2204), .B(n2582), .O(n1832));
  andx g1734(.A(n2208), .B(pi05), .O(n1833));
  andx g1735(.A(n2354), .B(n2436), .O(n1834));
  andx g1736(.A(pi00), .B(n2360), .O(n1835));
  andx g1737(.A(n2211), .B(n2210), .O(n1836));
  andx g1738(.A(n2213), .B(n2212), .O(n1837));
  andx g1739(.A(n2215), .B(n2214), .O(n1838));
  andx g1740(.A(n2217), .B(n2216), .O(n1839));
  andx g1741(.A(n2209), .B(n2335), .O(n1840));
  andx g1742(.A(n1557), .B(pi06), .O(n1841));
  andx g1743(.A(n2359), .B(n2438), .O(n1842));
  andx g1744(.A(pi00), .B(n2344), .O(n1843));
  andx g1745(.A(n2695), .B(n2521), .O(n1844));
  andx g1746(.A(n2218), .B(pi04), .O(n1845));
  andx g1747(.A(pi00), .B(n2764), .O(n1846));
  andx g1748(.A(pi02), .B(n2437), .O(n1847));
  andx g1749(.A(n2395), .B(n2439), .O(n1848));
  andx g1750(.A(pi00), .B(n2344), .O(n1849));
  andx g1751(.A(n2220), .B(n2523), .O(n1850));
  andx g1752(.A(n2221), .B(pi04), .O(n1851));
  andx g1753(.A(n2219), .B(n2478), .O(n1852));
  andx g1754(.A(n2222), .B(pi03), .O(n1853));
  andx g1755(.A(n2715), .B(n2523), .O(n1854));
  andx g1756(.A(pi04), .B(n2047), .O(n1855));
  andx g1757(.A(n2714), .B(pi04), .O(n1856));
  andx g1758(.A(n2065), .B(n2522), .O(n1857));
  andx g1759(.A(n2224), .B(n2476), .O(n1858));
  andx g1760(.A(n2225), .B(pi03), .O(n1859));
  andx g1761(.A(n2223), .B(n2582), .O(n1860));
  andx g1762(.A(n2226), .B(pi05), .O(n1861));
  andx g1763(.A(n2229), .B(n2228), .O(n1862));
  andx g1764(.A(n2231), .B(n2230), .O(n1863));
  andx g1765(.A(n2233), .B(n2232), .O(n1864));
  andx g1766(.A(n2227), .B(n2362), .O(n1865));
  andx g1767(.A(n1559), .B(pi06), .O(n1866));
  andx g1768(.A(n2382), .B(pi03), .O(n1867));
  andx g1769(.A(n1494), .B(n2478), .O(n1868));
  andx g1770(.A(n2150), .B(pi03), .O(n1869));
  andx g1771(.A(n2189), .B(n2477), .O(n1870));
  andx g1772(.A(n2234), .B(n2524), .O(n1871));
  andx g1773(.A(n2235), .B(pi04), .O(n1872));
  andx g1774(.A(n2075), .B(n2477), .O(n1873));
  andx g1775(.A(n2119), .B(pi03), .O(n1874));
  andx g1776(.A(n2706), .B(pi04), .O(n1875));
  andx g1777(.A(n2237), .B(n2522), .O(n1876));
  andx g1778(.A(n2236), .B(n2579), .O(n1877));
  andx g1779(.A(n2238), .B(pi05), .O(n1878));
  andx g1780(.A(n2241), .B(n2240), .O(n1879));
  orx  g1781(.A(pi03), .B(pi00), .O(n1880));
  andx g1782(.A(n2243), .B(n2242), .O(n1881));
  andx g1783(.A(n2245), .B(n2244), .O(n1882));
  andx g1784(.A(n2239), .B(n2353), .O(n1883));
  andx g1785(.A(n1561), .B(pi06), .O(n1884));
  andx g1786(.A(pi06), .B(pi01), .O(n1885));
  andx g1787(.A(n2332), .B(n2350), .O(n1886));
  andx g1788(.A(pi00), .B(n2331), .O(n1887));
  andx g1789(.A(pi06), .B(n2435), .O(n1888));
  andx g1790(.A(n1511), .B(n2680), .O(n1889));
  andx g1791(.A(n1516), .B(n2246), .O(n1890));
  andx g1792(.A(n2051), .B(n2335), .O(n1891));
  andx g1793(.A(pi06), .B(n2686), .O(n1892));
  andx g1794(.A(n2247), .B(n2479), .O(n1893));
  andx g1795(.A(n2248), .B(pi03), .O(n1894));
  andx g1796(.A(n1512), .B(pi06), .O(n1895));
  andx g1797(.A(n2167), .B(n2352), .O(n1896));
  andx g1798(.A(pi06), .B(n2389), .O(n1897));
  andx g1799(.A(n2341), .B(n2363), .O(n1898));
  andx g1800(.A(n2250), .B(n2480), .O(n1899));
  andx g1801(.A(n2251), .B(pi03), .O(n1900));
  andx g1802(.A(n2249), .B(n2524), .O(n1901));
  andx g1803(.A(n2252), .B(pi04), .O(n1902));
  andx g1804(.A(n2333), .B(n2439), .O(n1903));
  andx g1805(.A(pi00), .B(n2383), .O(n1904));
  andx g1806(.A(n2255), .B(n2254), .O(n1905));
  andx g1807(.A(pi01), .B(n2473), .O(n1906));
  andx g1808(.A(pi03), .B(n2355), .O(n1907));
  andx g1809(.A(n2257), .B(n2256), .O(n1908));
  andx g1810(.A(n2259), .B(n2258), .O(n1909));
  andx g1811(.A(n2253), .B(n2582), .O(n1910));
  andx g1812(.A(n1564), .B(pi05), .O(n1911));
  andx g1813(.A(pi01), .B(n2437), .O(n1912));
  andx g1814(.A(pi00), .B(n2384), .O(n1913));
  andx g1815(.A(n2704), .B(pi05), .O(n1914));
  andx g1816(.A(n1566), .B(n2583), .O(n1915));
  andx g1817(.A(n2066), .B(n2480), .O(n1916));
  andx g1818(.A(n2260), .B(pi03), .O(n1917));
  andx g1819(.A(pi00), .B(n2357), .O(n1918));
  andx g1820(.A(n2373), .B(n2432), .O(n1919));
  andx g1821(.A(n2136), .B(pi05), .O(n1920));
  andx g1822(.A(n2262), .B(n2580), .O(n1921));
  andx g1823(.A(n2381), .B(pi05), .O(n1922));
  andx g1824(.A(n2340), .B(n2576), .O(n1923));
  andx g1825(.A(n2263), .B(n2480), .O(n1924));
  andx g1826(.A(n2264), .B(pi03), .O(n1925));
  andx g1827(.A(n2261), .B(n2521), .O(n1926));
  andx g1828(.A(n2265), .B(pi04), .O(n1927));
  orx  g1829(.A(pi04), .B(pi03), .O(n1928));
  andx g1830(.A(n2268), .B(n2267), .O(n1929));
  andx g1831(.A(n2270), .B(n2269), .O(n1930));
  andx g1832(.A(n2272), .B(n2271), .O(n1931));
  andx g1833(.A(n2274), .B(n2273), .O(n1932));
  andx g1834(.A(n2266), .B(n2747), .O(n1933));
  andx g1835(.A(n1567), .B(pi06), .O(n1934));
  andx g1836(.A(n1514), .B(pi06), .O(n1935));
  andx g1837(.A(n2713), .B(n2350), .O(n1936));
  andx g1838(.A(n2705), .B(n2351), .O(n1937));
  andx g1839(.A(n2193), .B(pi06), .O(n1938));
  andx g1840(.A(n2275), .B(n2480), .O(n1939));
  andx g1841(.A(n2276), .B(pi03), .O(n1940));
  andx g1842(.A(n2703), .B(n2336), .O(n1941));
  andx g1843(.A(n1555), .B(pi06), .O(n1942));
  andx g1844(.A(n2251), .B(pi03), .O(n1943));
  andx g1845(.A(n2278), .B(n2478), .O(n1944));
  andx g1846(.A(n2277), .B(n2525), .O(n1945));
  andx g1847(.A(n2279), .B(pi04), .O(n1946));
  andx g1848(.A(n2282), .B(n2281), .O(n1947));
  andx g1849(.A(pi00), .B(n2343), .O(n1948));
  andx g1850(.A(n2342), .B(n2438), .O(n1949));
  andx g1851(.A(n2284), .B(n2283), .O(n1950));
  andx g1852(.A(n2286), .B(n2285), .O(n1951));
  andx g1853(.A(n2280), .B(n2583), .O(n1952));
  andx g1854(.A(n1569), .B(pi05), .O(n1953));
  andx g1855(.A(pi00), .B(n2358), .O(n1954));
  andx g1856(.A(n2379), .B(n2439), .O(n1955));
  andx g1857(.A(n1519), .B(pi03), .O(n1956));
  andx g1858(.A(n2287), .B(n2481), .O(n1957));
  andx g1859(.A(n2288), .B(n2523), .O(n1958));
  andx g1860(.A(n1571), .B(pi04), .O(n1959));
  andx g1861(.A(n2484), .B(n2436), .O(n1960));
  andx g1862(.A(pi03), .B(n2046), .O(n1961));
  andx g1863(.A(n2393), .B(n2439), .O(n1962));
  andx g1864(.A(n2382), .B(pi00), .O(n1963));
  andx g1865(.A(n2697), .B(pi03), .O(n1964));
  andx g1866(.A(n2291), .B(n2481), .O(n1965));
  andx g1867(.A(n2290), .B(n2525), .O(n1966));
  andx g1868(.A(n2292), .B(pi04), .O(n1967));
  andx g1869(.A(n2289), .B(n2581), .O(n1968));
  andx g1870(.A(n2293), .B(pi05), .O(n1969));
  andx g1871(.A(n2296), .B(n2295), .O(n1970));
  andx g1872(.A(n2298), .B(n2297), .O(n1971));
  andx g1873(.A(n2294), .B(n2331), .O(n1972));
  andx g1874(.A(n1572), .B(pi06), .O(n1973));
  andx g1875(.A(n2051), .B(pi04), .O(n1974));
  andx g1876(.A(n1512), .B(n2523), .O(n1975));
  andx g1877(.A(n2687), .B(n2526), .O(n1976));
  andx g1878(.A(n1517), .B(pi04), .O(n1977));
  andx g1879(.A(n2299), .B(n2481), .O(n1978));
  andx g1880(.A(n2300), .B(pi03), .O(n1979));
  andx g1881(.A(n2723), .B(pi04), .O(n1980));
  andx g1882(.A(n2092), .B(n2504), .O(n1981));
  andx g1883(.A(pi01), .B(n2526), .O(n1982));
  andx g1884(.A(n2381), .B(pi04), .O(n1983));
  andx g1885(.A(n2302), .B(n2479), .O(n1984));
  andx g1886(.A(n2303), .B(pi03), .O(n1985));
  andx g1887(.A(n2301), .B(n2583), .O(n1986));
  andx g1888(.A(n2304), .B(pi05), .O(n1987));
  andx g1889(.A(n2307), .B(n2306), .O(n1988));
  orx  g1890(.A(n1494), .B(pi04), .O(n1989));
  andx g1891(.A(n2309), .B(n2308), .O(n1990));
  andx g1892(.A(n2305), .B(n2336), .O(n1991));
  andx g1893(.A(n1574), .B(pi06), .O(n1992));
  andx g1894(.A(n1503), .B(n2524), .O(n1993));
  andx g1895(.A(n2092), .B(pi04), .O(n1994));
  andx g1896(.A(n2691), .B(n2526), .O(n1995));
  andx g1897(.A(n2262), .B(pi04), .O(n1996));
  andx g1898(.A(n2310), .B(n2481), .O(n1997));
  andx g1899(.A(n2311), .B(pi03), .O(n1998));
  andx g1900(.A(n1524), .B(n2524), .O(n1999));
  andx g1901(.A(n1550), .B(pi04), .O(n2000));
  andx g1902(.A(pi02), .B(n2526), .O(n2001));
  andx g1903(.A(pi04), .B(n2344), .O(n2002));
  andx g1904(.A(n2313), .B(n2476), .O(n2003));
  andx g1905(.A(n2314), .B(pi03), .O(n2004));
  andx g1906(.A(n2312), .B(n2583), .O(n2005));
  andx g1907(.A(n2315), .B(pi05), .O(n2006));
  andx g1908(.A(pi03), .B(n2521), .O(n2007));
  andx g1909(.A(pi04), .B(n2482), .O(n2008));
  andx g1910(.A(pi03), .B(n2388), .O(n2009));
  andx g1911(.A(n2341), .B(n2478), .O(n2010));
  andx g1912(.A(n2316), .B(n2353), .O(n2011));
  andx g1913(.A(n1577), .B(pi06), .O(n2012));
  andx g1914(.A(n1524), .B(pi04), .O(n2013));
  andx g1915(.A(n1579), .B(n2527), .O(n2014));
  andx g1916(.A(pi04), .B(n2703), .O(n2015));
  andx g1917(.A(n2092), .B(n2525), .O(n2016));
  andx g1918(.A(n2317), .B(n2482), .O(n2017));
  andx g1919(.A(n2318), .B(pi03), .O(n2018));
  andx g1920(.A(n2687), .B(pi04), .O(n2019));
  andx g1921(.A(n2707), .B(n2520), .O(n2020));
  andx g1922(.A(n2320), .B(n2479), .O(n2021));
  andx g1923(.A(n2069), .B(pi03), .O(n2022));
  andx g1924(.A(n2319), .B(n2582), .O(n2023));
  andx g1925(.A(n2321), .B(pi05), .O(n2024));
  andx g1926(.A(n2322), .B(n2362), .O(n2025));
  andx g1927(.A(n1580), .B(pi06), .O(n2026));
  andx g1928(.A(n1524), .B(pi03), .O(n2027));
  andx g1929(.A(n1535), .B(n2482), .O(n2028));
  andx g1930(.A(n1491), .B(pi03), .O(n2029));
  andx g1931(.A(n2707), .B(n2479), .O(n2030));
  andx g1932(.A(n2323), .B(n2525), .O(n2031));
  andx g1933(.A(n2324), .B(pi04), .O(n2032));
  andx g1934(.A(n2325), .B(n2584), .O(n2033));
  andx g1935(.A(n1582), .B(pi05), .O(n2034));
  andx g1936(.A(n2326), .B(n2331), .O(n2035));
  andx g1937(.A(n1583), .B(pi06), .O(n2036));
  andx g1938(.A(n2328), .B(n2327), .O(n2037));
  orx  g1939(.A(pi05), .B(n1510), .O(n2038));
  andx g1940(.A(n2072), .B(n2362), .O(n2039));
  andx g1941(.A(n2683), .B(pi06), .O(n2040));
  andx g1942(.A(n2683), .B(pi06), .O(n2041));
  andx g1943(.A(n2073), .B(n2352), .O(n2042));
  andx g1944(.A(n2683), .B(pi06), .O(n2043));
  andx g1945(.A(n2074), .B(n2349), .O(n2044));
  orx  g1946(.A(pi00), .B(n2344), .O(n2045));
  orx  g1947(.A(n2390), .B(n2710), .O(n2046));
  orx  g1948(.A(pi00), .B(n2760), .O(n2047));
  orx  g1949(.A(n2385), .B(n2443), .O(n2048));
  orx  g1950(.A(n2382), .B(n2443), .O(n2049));
  orx  g1951(.A(n2389), .B(n2443), .O(n2050));
  orx  g1952(.A(n2342), .B(n2443), .O(n2051));
  orx  g1953(.A(n2710), .B(n2366), .O(n2052));
  orx  g1954(.A(n2341), .B(n2719), .O(n2053));
  orx  g1955(.A(n2693), .B(n2530), .O(n2054));
  orx  g1956(.A(n2392), .B(n2444), .O(n2055));
  orx  g1957(.A(pi01), .B(n2444), .O(n2056));
  orx  g1958(.A(n2709), .B(n1488), .O(n2057));
  orx  g1959(.A(n2719), .B(n2333), .O(n2058));
  orx  g1960(.A(n1540), .B(n1490), .O(n2059));
  orx  g1961(.A(n1493), .B(n1492), .O(n2060));
  orx  g1962(.A(n2706), .B(n2530), .O(n2061));
  orx  g1963(.A(n1514), .B(n2530), .O(n2062));
  orx  g1964(.A(n1494), .B(n2530), .O(n2063));
  orx  g1965(.A(n1555), .B(pi04), .O(n2064));
  orx  g1966(.A(n2340), .B(n2701), .O(n2065));
  orx  g1967(.A(n1495), .B(n2707), .O(n2066));
  orx  g1968(.A(n2709), .B(n2485), .O(n2067));
  orx  g1969(.A(n1518), .B(n1576), .O(n2068));
  orx  g1970(.A(n2342), .B(n2531), .O(n2069));
  orx  g1971(.A(n1506), .B(n2388), .O(n2070));
  orx  g1972(.A(n1496), .B(n2531), .O(n2071));
  orx  g1973(.A(n1498), .B(pi05), .O(n2072));
  orx  g1974(.A(n1499), .B(pi03), .O(n2073));
  orx  g1975(.A(n1499), .B(n1497), .O(n2074));
  orx  g1976(.A(n1592), .B(n1593), .O(n2075));
  orx  g1977(.A(n1594), .B(n1595), .O(n2076));
  orx  g1978(.A(n1596), .B(n1597), .O(n2077));
  orx  g1979(.A(n1598), .B(n1599), .O(n2078));
  orx  g1980(.A(n1602), .B(n1603), .O(n2079));
  orx  g1981(.A(n1604), .B(n1605), .O(n2080));
  orx  g1982(.A(n1606), .B(n1607), .O(n2081));
  orx  g1983(.A(n1608), .B(n1609), .O(n2082));
  orx  g1984(.A(n1610), .B(n1611), .O(n2083));
  orx  g1985(.A(n1612), .B(n1613), .O(n2084));
  orx  g1986(.A(pi04), .B(n2715), .O(n2085));
  orx  g1987(.A(n2499), .B(n1519), .O(n2086));
  orx  g1988(.A(pi01), .B(n2444), .O(n2087));
  orx  g1989(.A(pi00), .B(n2381), .O(n2088));
  orx  g1990(.A(pi03), .B(n1616), .O(n2089));
  orx  g1991(.A(n2458), .B(n1520), .O(n2090));
  orx  g1992(.A(n1621), .B(n1622), .O(n2091));
  orx  g1993(.A(n1623), .B(n1624), .O(n2092));
  orx  g1994(.A(n1627), .B(n1628), .O(n2093));
  orx  g1995(.A(n1629), .B(n1630), .O(n2094));
  orx  g1996(.A(n1631), .B(n1632), .O(n2095));
  orx  g1997(.A(n1633), .B(n1634), .O(n2096));
  orx  g1998(.A(n1637), .B(n1638), .O(n2097));
  orx  g1999(.A(n1639), .B(n1640), .O(n2098));
  orx  g2000(.A(n1641), .B(n1642), .O(n2099));
  orx  g2001(.A(n2499), .B(n1643), .O(n2100));
  orx  g2002(.A(pi04), .B(n2724), .O(n2101));
  orx  g2003(.A(pi04), .B(n2717), .O(n2102));
  orx  g2004(.A(n2687), .B(n2531), .O(n2103));
  orx  g2005(.A(pi03), .B(n1644), .O(n2104));
  orx  g2006(.A(n2457), .B(n1645), .O(n2105));
  orx  g2007(.A(n1649), .B(n1650), .O(n2106));
  orx  g2008(.A(n1651), .B(n1652), .O(n2107));
  orx  g2009(.A(n1653), .B(n1654), .O(n2108));
  orx  g2010(.A(n1657), .B(n1658), .O(n2109));
  orx  g2011(.A(n1659), .B(n1660), .O(n2110));
  orx  g2012(.A(n1661), .B(n1662), .O(n2111));
  orx  g2013(.A(n1663), .B(n1664), .O(n2112));
  orx  g2014(.A(n1665), .B(n1666), .O(n2113));
  orx  g2015(.A(n1667), .B(n1668), .O(n2114));
  orx  g2016(.A(pi04), .B(n1524), .O(n2115));
  orx  g2017(.A(n2499), .B(n1512), .O(n2116));
  orx  g2018(.A(pi03), .B(n1671), .O(n2117));
  orx  g2019(.A(n2457), .B(n1527), .O(n2118));
  orx  g2020(.A(n1675), .B(n1676), .O(n2119));
  orx  g2021(.A(n1677), .B(n1678), .O(n2120));
  orx  g2022(.A(n1679), .B(n1680), .O(n2121));
  orx  g2023(.A(n1681), .B(n1682), .O(n2122));
  orx  g2024(.A(n1683), .B(n1684), .O(n2123));
  orx  g2025(.A(n1685), .B(n1686), .O(n2124));
  orx  g2026(.A(n1687), .B(n1688), .O(n2125));
  orx  g2027(.A(n1689), .B(n1690), .O(n2126));
  orx  g2028(.A(n2404), .B(n2384), .O(n2127));
  orx  g2029(.A(pi00), .B(n2365), .O(n2128));
  orx  g2030(.A(n1692), .B(n1693), .O(n2129));
  orx  g2031(.A(n1694), .B(n1695), .O(n2130));
  orx  g2032(.A(n1696), .B(n1697), .O(n2131));
  orx  g2033(.A(n2457), .B(n1700), .O(n2132));
  orx  g2034(.A(pi03), .B(n1530), .O(n2133));
  orx  g2035(.A(pi04), .B(n1701), .O(n2134));
  orx  g2036(.A(n2698), .B(n2531), .O(n2135));
  orx  g2037(.A(n1705), .B(n1706), .O(n2136));
  orx  g2038(.A(n1708), .B(n1707), .O(n2137));
  orx  g2039(.A(n1709), .B(n1710), .O(n2138));
  orx  g2040(.A(n1714), .B(n1713), .O(n2139));
  orx  g2041(.A(n1715), .B(n1716), .O(n2140));
  orx  g2042(.A(n1717), .B(n1718), .O(n2141));
  orx  g2043(.A(n1719), .B(n1720), .O(n2142));
  orx  g2044(.A(n1721), .B(n1722), .O(n2143));
  orx  g2045(.A(pi02), .B(n2486), .O(n2144));
  orx  g2046(.A(pi03), .B(n2382), .O(n2145));
  orx  g2047(.A(n2403), .B(n2531), .O(n2146));
  orx  g2048(.A(pi04), .B(n1723), .O(n2147));
  orx  g2049(.A(n1533), .B(n2332), .O(n2148));
  orx  g2050(.A(n1724), .B(n2678), .O(n2149));
  orx  g2051(.A(n1730), .B(n1731), .O(n2150));
  orx  g2052(.A(n1734), .B(n1735), .O(n2151));
  orx  g2053(.A(n1736), .B(n1737), .O(n2152));
  orx  g2054(.A(n1738), .B(n1739), .O(n2153));
  orx  g2055(.A(n1740), .B(n1741), .O(n2154));
  orx  g2056(.A(n1742), .B(n1743), .O(n2155));
  orx  g2057(.A(n1744), .B(n1745), .O(n2156));
  orx  g2058(.A(n1746), .B(n1747), .O(n2157));
  orx  g2059(.A(pi04), .B(n2586), .O(n2158));
  orx  g2060(.A(n2498), .B(n1508), .O(n2159));
  orx  g2061(.A(pi03), .B(n2365), .O(n2160));
  orx  g2062(.A(n2712), .B(n2486), .O(n2161));
  orx  g2063(.A(pi00), .B(n2532), .O(n2162));
  orx  g2064(.A(pi04), .B(n1749), .O(n2163));
  orx  g2065(.A(n1753), .B(n1754), .O(n2164));
  orx  g2066(.A(n1757), .B(n1758), .O(n2165));
  orx  g2067(.A(n1759), .B(n1760), .O(n2166));
  orx  g2068(.A(n1763), .B(n1764), .O(n2167));
  orx  g2069(.A(n1765), .B(n1766), .O(n2168));
  orx  g2070(.A(n1767), .B(n1768), .O(n2169));
  orx  g2071(.A(n1769), .B(n1770), .O(n2170));
  orx  g2072(.A(pi04), .B(n1491), .O(n2171));
  orx  g2073(.A(n2498), .B(n1771), .O(n2172));
  orx  g2074(.A(pi04), .B(n1535), .O(n2173));
  orx  g2075(.A(n2498), .B(n2686), .O(n2174));
  orx  g2076(.A(pi03), .B(n1772), .O(n2175));
  orx  g2077(.A(n2757), .B(n1773), .O(n2176));
  orx  g2078(.A(n1779), .B(n1780), .O(n2177));
  orx  g2079(.A(n1781), .B(n1782), .O(n2178));
  orx  g2080(.A(n1783), .B(n1784), .O(n2179));
  orx  g2081(.A(n1785), .B(n1786), .O(n2180));
  orx  g2082(.A(n1787), .B(n1788), .O(n2181));
  orx  g2083(.A(pi00), .B(n2393), .O(n2182));
  orx  g2084(.A(n2380), .B(n2444), .O(n2183));
  orx  g2085(.A(n2497), .B(n2686), .O(n2184));
  orx  g2086(.A(pi04), .B(n1544), .O(n2185));
  orx  g2087(.A(pi03), .B(n1545), .O(n2186));
  orx  g2088(.A(n2476), .B(n1790), .O(n2187));
  orx  g2089(.A(n1794), .B(n1795), .O(n2188));
  orx  g2090(.A(n1796), .B(n1797), .O(n2189));
  orx  g2091(.A(n1798), .B(n1799), .O(n2190));
  orx  g2092(.A(n1800), .B(n1801), .O(n2191));
  orx  g2093(.A(n1802), .B(n1803), .O(n2192));
  orx  g2094(.A(n1804), .B(n1805), .O(n2193));
  orx  g2095(.A(n1806), .B(n1807), .O(n2194));
  orx  g2096(.A(n1808), .B(n1809), .O(n2195));
  orx  g2097(.A(n1810), .B(n1811), .O(n2196));
  orx  g2098(.A(pi03), .B(n1547), .O(n2197));
  orx  g2099(.A(n2467), .B(n1550), .O(n2198));
  orx  g2100(.A(n2687), .B(n2757), .O(n2199));
  orx  g2101(.A(pi03), .B(n1530), .O(n2200));
  orx  g2102(.A(pi04), .B(n1814), .O(n2201));
  orx  g2103(.A(n2497), .B(n1815), .O(n2202));
  orx  g2104(.A(n2016), .B(n1819), .O(n2203));
  orx  g2105(.A(n1820), .B(n1821), .O(n2204));
  orx  g2106(.A(n1824), .B(n1825), .O(n2205));
  orx  g2107(.A(n1826), .B(n1827), .O(n2206));
  orx  g2108(.A(n1828), .B(n1829), .O(n2207));
  orx  g2109(.A(n1830), .B(n1831), .O(n2208));
  orx  g2110(.A(n1832), .B(n1833), .O(n2209));
  orx  g2111(.A(pi04), .B(n2721), .O(n2210));
  orx  g2112(.A(n2497), .B(n1554), .O(n2211));
  orx  g2113(.A(n2357), .B(n2444), .O(n2212));
  orx  g2114(.A(pi00), .B(n2360), .O(n2213));
  orx  g2115(.A(n2497), .B(n2390), .O(n2214));
  orx  g2116(.A(pi04), .B(n1837), .O(n2215));
  orx  g2117(.A(pi03), .B(n1836), .O(n2216));
  orx  g2118(.A(n2456), .B(n1838), .O(n2217));
  orx  g2119(.A(n1842), .B(n1843), .O(n2218));
  orx  g2120(.A(n1844), .B(n1845), .O(n2219));
  orx  g2121(.A(n1846), .B(n1847), .O(n2220));
  orx  g2122(.A(n1848), .B(n1849), .O(n2221));
  orx  g2123(.A(n1850), .B(n1851), .O(n2222));
  orx  g2124(.A(n1852), .B(n1853), .O(n2223));
  orx  g2125(.A(n1854), .B(n1855), .O(n2224));
  orx  g2126(.A(n1856), .B(n1857), .O(n2225));
  orx  g2127(.A(n1858), .B(n1859), .O(n2226));
  orx  g2128(.A(n1860), .B(n1861), .O(n2227));
  orx  g2129(.A(pi04), .B(n2706), .O(n2228));
  orx  g2130(.A(n2341), .B(n2532), .O(n2229));
  orx  g2131(.A(pi04), .B(n2723), .O(n2230));
  orx  g2132(.A(n2495), .B(n2686), .O(n2231));
  orx  g2133(.A(pi03), .B(n1862), .O(n2232));
  orx  g2134(.A(n2456), .B(n1863), .O(n2233));
  orx  g2135(.A(n1867), .B(n1868), .O(n2234));
  orx  g2136(.A(n1869), .B(n1870), .O(n2235));
  orx  g2137(.A(n1871), .B(n1872), .O(n2236));
  orx  g2138(.A(n1873), .B(n1874), .O(n2237));
  orx  g2139(.A(n1875), .B(n1876), .O(n2238));
  orx  g2140(.A(n1877), .B(n1878), .O(n2239));
  orx  g2141(.A(n2456), .B(n1700), .O(n2240));
  orx  g2142(.A(pi03), .B(n2720), .O(n2241));
  orx  g2143(.A(n2388), .B(n2728), .O(n2242));
  orx  g2144(.A(n2340), .B(n1880), .O(n2243));
  orx  g2145(.A(pi04), .B(n1879), .O(n2244));
  orx  g2146(.A(n2496), .B(n1881), .O(n2245));
  orx  g2147(.A(n1885), .B(n1886), .O(n2246));
  orx  g2148(.A(n1889), .B(n1890), .O(n2247));
  orx  g2149(.A(n1892), .B(n1891), .O(n2248));
  orx  g2150(.A(n1893), .B(n1894), .O(n2249));
  orx  g2151(.A(n1895), .B(n1896), .O(n2250));
  orx  g2152(.A(n1897), .B(n1898), .O(n2251));
  orx  g2153(.A(n1899), .B(n1900), .O(n2252));
  orx  g2154(.A(n1901), .B(n1902), .O(n2253));
  orx  g2155(.A(n2456), .B(n1554), .O(n2254));
  orx  g2156(.A(pi03), .B(n1563), .O(n2255));
  orx  g2157(.A(pi00), .B(n2366), .O(n2256));
  orx  g2158(.A(n2403), .B(n1515), .O(n2257));
  orx  g2159(.A(pi04), .B(n1905), .O(n2258));
  orx  g2160(.A(n2496), .B(n1908), .O(n2259));
  orx  g2161(.A(n1914), .B(n1915), .O(n2260));
  orx  g2162(.A(n1916), .B(n1917), .O(n2261));
  orx  g2163(.A(n1918), .B(n1919), .O(n2262));
  orx  g2164(.A(n1920), .B(n1921), .O(n2263));
  orx  g2165(.A(n1922), .B(n1923), .O(n2264));
  orx  g2166(.A(n1924), .B(n1925), .O(n2265));
  orx  g2167(.A(n1926), .B(n1927), .O(n2266));
  orx  g2168(.A(n2541), .B(n2676), .O(n2267));
  orx  g2169(.A(n1509), .B(n1928), .O(n2268));
  orx  g2170(.A(pi03), .B(n2381), .O(n2269));
  orx  g2171(.A(n2455), .B(n1514), .O(n2270));
  orx  g2172(.A(n2455), .B(n2389), .O(n2271));
  orx  g2173(.A(pi03), .B(n2700), .O(n2272));
  orx  g2174(.A(pi04), .B(n1930), .O(n2273));
  orx  g2175(.A(n2496), .B(n1931), .O(n2274));
  orx  g2176(.A(n1935), .B(n1936), .O(n2275));
  orx  g2177(.A(n1938), .B(n1937), .O(n2276));
  orx  g2178(.A(n1939), .B(n1940), .O(n2277));
  orx  g2179(.A(n1942), .B(n1941), .O(n2278));
  orx  g2180(.A(n1943), .B(n1944), .O(n2279));
  orx  g2181(.A(n1945), .B(n1946), .O(n2280));
  orx  g2182(.A(n2455), .B(n1501), .O(n2281));
  orx  g2183(.A(pi03), .B(n2343), .O(n2282));
  orx  g2184(.A(pi03), .B(n1563), .O(n2283));
  orx  g2185(.A(n2455), .B(n1517), .O(n2284));
  orx  g2186(.A(pi04), .B(n1947), .O(n2285));
  orx  g2187(.A(n2495), .B(n1950), .O(n2286));
  orx  g2188(.A(n1954), .B(n1955), .O(n2287));
  orx  g2189(.A(n1956), .B(n1957), .O(n2288));
  orx  g2190(.A(n1958), .B(n1959), .O(n2289));
  orx  g2191(.A(n1960), .B(n1961), .O(n2290));
  orx  g2192(.A(n1962), .B(n1963), .O(n2291));
  orx  g2193(.A(n1964), .B(n1965), .O(n2292));
  orx  g2194(.A(n1966), .B(n1967), .O(n2293));
  orx  g2195(.A(n1968), .B(n1969), .O(n2294));
  orx  g2196(.A(pi03), .B(n2716), .O(n2295));
  orx  g2197(.A(n2454), .B(n2692), .O(n2296));
  orx  g2198(.A(pi04), .B(n1970), .O(n2297));
  orx  g2199(.A(n1496), .B(n2532), .O(n2298));
  orx  g2200(.A(n1974), .B(n1975), .O(n2299));
  orx  g2201(.A(n1976), .B(n1977), .O(n2300));
  orx  g2202(.A(n1978), .B(n1979), .O(n2301));
  orx  g2203(.A(n1980), .B(n1981), .O(n2302));
  orx  g2204(.A(n1982), .B(n1983), .O(n2303));
  orx  g2205(.A(n1984), .B(n1985), .O(n2304));
  orx  g2206(.A(n1986), .B(n1987), .O(n2305));
  orx  g2207(.A(pi02), .B(pi04), .O(n2306));
  orx  g2208(.A(n2495), .B(n2388), .O(n2307));
  orx  g2209(.A(pi03), .B(n1989), .O(n2308));
  orx  g2210(.A(n2454), .B(n1988), .O(n2309));
  orx  g2211(.A(n1993), .B(n1994), .O(n2310));
  orx  g2212(.A(n1995), .B(n1996), .O(n2311));
  orx  g2213(.A(n1997), .B(n1998), .O(n2312));
  orx  g2214(.A(n1999), .B(n2000), .O(n2313));
  orx  g2215(.A(n2001), .B(n2002), .O(n2314));
  orx  g2216(.A(n2003), .B(n2004), .O(n2315));
  orx  g2217(.A(n2005), .B(n2006), .O(n2316));
  orx  g2218(.A(n2013), .B(n2014), .O(n2317));
  orx  g2219(.A(n2015), .B(n2016), .O(n2318));
  orx  g2220(.A(n2017), .B(n2018), .O(n2319));
  orx  g2221(.A(n2019), .B(n2020), .O(n2320));
  orx  g2222(.A(n2021), .B(n2022), .O(n2321));
  orx  g2223(.A(n2023), .B(n2024), .O(n2322));
  orx  g2224(.A(n2027), .B(n2028), .O(n2323));
  orx  g2225(.A(n2029), .B(n2030), .O(n2324));
  orx  g2226(.A(n2031), .B(n2032), .O(n2325));
  orx  g2227(.A(n2033), .B(n2034), .O(n2326));
  orx  g2228(.A(pi04), .B(n2379), .O(n2327));
  orx  g2229(.A(n2495), .B(n2707), .O(n2328));
  invx g2230(.A(n2350), .O(n2329));
  invx g2231(.A(pi02), .O(n2330));
  invx g2232(.A(n2334), .O(n2331));
  invx g2233(.A(n2381), .O(n2332));
  invx g2234(.A(n1511), .O(n2333));
  invx g2235(.A(n2349), .O(n2334));
  invx g2236(.A(n2334), .O(n2335));
  invx g2237(.A(n2334), .O(n2336));
  invx g2238(.A(n2345), .O(n2337));
  invx g2239(.A(n2337), .O(n2338));
  invx g2240(.A(n2337), .O(n2339));
  invx g2241(.A(n2343), .O(n2340));
  invx g2242(.A(n1504), .O(n2341));
  invx g2243(.A(n1504), .O(n2342));
  invx g2244(.A(n2342), .O(n2343));
  invx g2245(.A(n2342), .O(n2344));
  invx g2246(.A(n181), .O(n2345));
  invx g2247(.A(n2345), .O(n2346));
  invx g2248(.A(n2345), .O(n2347));
  invx g2249(.A(n2345), .O(n2348));
  invx g2250(.A(pi06), .O(n2349));
  invx g2251(.A(pi06), .O(n2350));
  invx g2252(.A(n2334), .O(n2351));
  invx g2253(.A(n2329), .O(n2352));
  invx g2254(.A(n2334), .O(n2353));
  invx g2255(.A(pi01), .O(n2354));
  invx g2256(.A(pi01), .O(n2355));
  invx g2257(.A(pi01), .O(n2356));
  invx g2258(.A(pi01), .O(n2357));
  invx g2259(.A(pi02), .O(n2358));
  invx g2260(.A(pi02), .O(n2359));
  invx g2261(.A(pi02), .O(n2360));
  invx g2262(.A(pi02), .O(n2361));
  invx g2263(.A(pi06), .O(n2362));
  invx g2264(.A(pi06), .O(n2363));
  bufx g2265(.A(n2367), .O(n2364));
  bufx g2266(.A(n164), .O(n2365));
  bufx g2267(.A(n2718), .O(n2366));
  bufx g2268(.A(n2819), .O(n2367));
  bufx g2269(.A(n2396), .O(n2368));
  bufx g2270(.A(n2396), .O(n2369));
  bufx g2271(.A(n2727), .O(n2370));
  invx g2272(.A(n2365), .O(n2371));
  invx g2273(.A(n2371), .O(n2372));
  invx g2274(.A(n2371), .O(n2373));
  invx g2275(.A(n2399), .O(n2374));
  invx g2276(.A(n2399), .O(n2375));
  invx g2277(.A(n2399), .O(n2376));
  bufx g2278(.A(n2699), .O(n2377));
  bufx g2279(.A(n2699), .O(n2378));
  bufx g2280(.A(n1485), .O(n2379));
  bufx g2281(.A(n1485), .O(n2380));
  bufx g2282(.A(n1511), .O(n2381));
  bufx g2283(.A(n1511), .O(n2382));
  bufx g2284(.A(n2371), .O(n2383));
  bufx g2285(.A(n2371), .O(n2384));
  bufx g2286(.A(n2371), .O(n2385));
  bufx g2287(.A(n183), .O(n2386));
  bufx g2288(.A(n183), .O(n2387));
  bufx g2289(.A(n2688), .O(n2388));
  bufx g2290(.A(n2688), .O(n2389));
  bufx g2291(.A(n2688), .O(n2390));
  invx g2292(.A(n1484), .O(n2391));
  invx g2293(.A(n2391), .O(n2392));
  invx g2294(.A(n2391), .O(n2393));
  invx g2295(.A(n2391), .O(n2394));
  invx g2296(.A(n2391), .O(n2395));
  invx g2297(.A(n207), .O(n2396));
  invx g2298(.A(n2396), .O(n2397));
  invx g2299(.A(n2396), .O(n2398));
  invx g2300(.A(n2819), .O(n2399));
  invx g2301(.A(n2399), .O(n2400));
  invx g2302(.A(n2399), .O(n2401));
  invx g2303(.A(n2399), .O(n2402));
  invx g2304(.A(n2452), .O(n2403));
  invx g2305(.A(n2452), .O(n2404));
  invx g2306(.A(n2452), .O(n2405));
  invx g2307(.A(n2451), .O(n2406));
  invx g2308(.A(n2451), .O(n2407));
  invx g2309(.A(n2451), .O(n2408));
  invx g2310(.A(n2445), .O(n2409));
  invx g2311(.A(n2449), .O(n2410));
  invx g2312(.A(n2450), .O(n2411));
  invx g2313(.A(n2451), .O(n2412));
  invx g2314(.A(n2446), .O(n2413));
  invx g2315(.A(n2450), .O(n2414));
  invx g2316(.A(n2450), .O(n2415));
  invx g2317(.A(n2450), .O(n2416));
  invx g2318(.A(n2449), .O(n2417));
  invx g2319(.A(n2449), .O(n2418));
  invx g2320(.A(n2449), .O(n2419));
  invx g2321(.A(n2445), .O(n2420));
  invx g2322(.A(n2447), .O(n2421));
  invx g2323(.A(n2449), .O(n2422));
  invx g2324(.A(n2448), .O(n2423));
  invx g2325(.A(n2448), .O(n2424));
  invx g2326(.A(n2448), .O(n2425));
  invx g2327(.A(n2447), .O(n2426));
  invx g2328(.A(n2446), .O(n2427));
  invx g2329(.A(n2448), .O(n2428));
  invx g2330(.A(n2451), .O(n2429));
  invx g2331(.A(n2445), .O(n2430));
  invx g2332(.A(n2447), .O(n2431));
  invx g2333(.A(n2447), .O(n2432));
  invx g2334(.A(n2447), .O(n2433));
  invx g2335(.A(n2446), .O(n2434));
  invx g2336(.A(n2446), .O(n2435));
  invx g2337(.A(n2446), .O(n2436));
  invx g2338(.A(n2446), .O(n2437));
  invx g2339(.A(n2448), .O(n2438));
  invx g2340(.A(n2450), .O(n2439));
  invx g2341(.A(n2451), .O(n2440));
  invx g2342(.A(n2452), .O(n2441));
  invx g2343(.A(n2452), .O(n2442));
  invx g2344(.A(n2445), .O(n2443));
  invx g2345(.A(n2445), .O(n2444));
  invx g2346(.A(n2453), .O(n2445));
  invx g2347(.A(n2429), .O(n2446));
  invx g2348(.A(n2430), .O(n2447));
  invx g2349(.A(n2420), .O(n2448));
  invx g2350(.A(n2453), .O(n2449));
  invx g2351(.A(n2453), .O(n2450));
  invx g2352(.A(n2765), .O(n2451));
  invx g2353(.A(n2765), .O(n2452));
  invx g2354(.A(n2452), .O(n2453));
  invx g2355(.A(n2493), .O(n2454));
  invx g2356(.A(n2493), .O(n2455));
  invx g2357(.A(n2493), .O(n2456));
  invx g2358(.A(n2492), .O(n2457));
  invx g2359(.A(n2492), .O(n2458));
  invx g2360(.A(n2492), .O(n2459));
  invx g2361(.A(n2488), .O(n2460));
  invx g2362(.A(n2493), .O(n2461));
  invx g2363(.A(n2489), .O(n2462));
  invx g2364(.A(n2490), .O(n2463));
  invx g2365(.A(n2491), .O(n2464));
  invx g2366(.A(n2493), .O(n2465));
  invx g2367(.A(n2489), .O(n2466));
  invx g2368(.A(n2490), .O(n2467));
  invx g2369(.A(n2491), .O(n2468));
  invx g2370(.A(n2491), .O(n2469));
  invx g2371(.A(n2491), .O(n2470));
  invx g2372(.A(n2490), .O(n2471));
  invx g2373(.A(n2490), .O(n2472));
  invx g2374(.A(n2490), .O(n2473));
  invx g2375(.A(n2489), .O(n2474));
  invx g2376(.A(n2489), .O(n2475));
  invx g2377(.A(n2489), .O(n2476));
  invx g2378(.A(n2491), .O(n2477));
  invx g2379(.A(n2492), .O(n2478));
  invx g2380(.A(n2488), .O(n2479));
  invx g2381(.A(n2488), .O(n2480));
  invx g2382(.A(n2488), .O(n2481));
  invx g2383(.A(n2488), .O(n2482));
  invx g2384(.A(n2487), .O(n2483));
  invx g2385(.A(n2492), .O(n2484));
  invx g2386(.A(n2487), .O(n2485));
  invx g2387(.A(n2487), .O(n2486));
  invx g2388(.A(n2757), .O(n2487));
  invx g2389(.A(n2484), .O(n2488));
  invx g2390(.A(n2494), .O(n2489));
  invx g2391(.A(n2494), .O(n2490));
  invx g2392(.A(n2494), .O(n2491));
  invx g2393(.A(n2483), .O(n2492));
  invx g2394(.A(n2494), .O(n2493));
  invx g2395(.A(n2487), .O(n2494));
  invx g2396(.A(n2537), .O(n2495));
  invx g2397(.A(n2539), .O(n2496));
  invx g2398(.A(n2539), .O(n2497));
  invx g2399(.A(n2539), .O(n2498));
  invx g2400(.A(n2539), .O(n2499));
  invx g2401(.A(n2534), .O(n2500));
  invx g2402(.A(n2534), .O(n2501));
  invx g2403(.A(n2533), .O(n2502));
  invx g2404(.A(n2538), .O(n2503));
  invx g2405(.A(n2538), .O(n2504));
  invx g2406(.A(n2538), .O(n2505));
  invx g2407(.A(n2537), .O(n2506));
  invx g2408(.A(n2534), .O(n2507));
  invx g2409(.A(n2537), .O(n2508));
  invx g2410(.A(n2537), .O(n2509));
  invx g2411(.A(n2537), .O(n2510));
  invx g2412(.A(n2536), .O(n2511));
  invx g2413(.A(n2536), .O(n2512));
  invx g2414(.A(n2536), .O(n2513));
  invx g2415(.A(n2535), .O(n2514));
  invx g2416(.A(n2535), .O(n2515));
  invx g2417(.A(n2535), .O(n2516));
  invx g2418(.A(n2534), .O(n2517));
  invx g2419(.A(n2534), .O(n2518));
  invx g2420(.A(n2534), .O(n2519));
  invx g2421(.A(n2533), .O(n2520));
  invx g2422(.A(n2538), .O(n2521));
  invx g2423(.A(n2539), .O(n2522));
  invx g2424(.A(n2537), .O(n2523));
  invx g2425(.A(n2533), .O(n2524));
  invx g2426(.A(n2533), .O(n2525));
  invx g2427(.A(n2533), .O(n2526));
  invx g2428(.A(n2538), .O(n2527));
  invx g2429(.A(n2535), .O(n2528));
  invx g2430(.A(n2536), .O(n2529));
  invx g2431(.A(n2535), .O(n2530));
  invx g2432(.A(n2536), .O(n2531));
  invx g2433(.A(n2533), .O(n2532));
  invx g2434(.A(n2751), .O(n2533));
  invx g2435(.A(n2540), .O(n2534));
  invx g2436(.A(n2540), .O(n2535));
  invx g2437(.A(n2540), .O(n2536));
  invx g2438(.A(n2540), .O(n2537));
  invx g2439(.A(n2520), .O(n2538));
  invx g2440(.A(n2751), .O(n2539));
  invx g2441(.A(n2539), .O(n2540));
  invx g2442(.A(n2588), .O(n2541));
  invx g2443(.A(n2587), .O(n2542));
  invx g2444(.A(n2593), .O(n2543));
  invx g2445(.A(n2596), .O(n2544));
  invx g2446(.A(n2596), .O(n2545));
  invx g2447(.A(n2596), .O(n2546));
  invx g2448(.A(n2595), .O(n2547));
  invx g2449(.A(n2595), .O(n2548));
  invx g2450(.A(n2595), .O(n2549));
  invx g2451(.A(n2594), .O(n2550));
  invx g2452(.A(n2594), .O(n2551));
  invx g2453(.A(n2594), .O(n2552));
  invx g2454(.A(n2591), .O(n2553));
  invx g2455(.A(n2591), .O(n2554));
  invx g2456(.A(n2592), .O(n2555));
  invx g2457(.A(n2593), .O(n2556));
  invx g2458(.A(n2593), .O(n2557));
  invx g2459(.A(n2593), .O(n2558));
  invx g2460(.A(n2592), .O(n2559));
  invx g2461(.A(n2592), .O(n2560));
  invx g2462(.A(n2592), .O(n2561));
  invx g2463(.A(n2591), .O(n2562));
  invx g2464(.A(n2591), .O(n2563));
  invx g2465(.A(n2591), .O(n2564));
  invx g2466(.A(n2589), .O(n2565));
  invx g2467(.A(n2590), .O(n2566));
  invx g2468(.A(n2590), .O(n2567));
  invx g2469(.A(n2590), .O(n2568));
  invx g2470(.A(n2590), .O(n2569));
  invx g2471(.A(n2589), .O(n2570));
  invx g2472(.A(n2589), .O(n2571));
  invx g2473(.A(n2589), .O(n2572));
  invx g2474(.A(n2596), .O(n2573));
  invx g2475(.A(n2595), .O(n2574));
  invx g2476(.A(n2588), .O(n2575));
  invx g2477(.A(n2588), .O(n2576));
  invx g2478(.A(n2588), .O(n2577));
  invx g2479(.A(n2588), .O(n2578));
  invx g2480(.A(n2587), .O(n2579));
  invx g2481(.A(n2587), .O(n2580));
  invx g2482(.A(n2587), .O(n2581));
  invx g2483(.A(n2593), .O(n2582));
  invx g2484(.A(n2594), .O(n2583));
  invx g2485(.A(n2587), .O(n2584));
  invx g2486(.A(n2595), .O(n2585));
  invx g2487(.A(n2592), .O(n2586));
  invx g2488(.A(n2744), .O(n2587));
  invx g2489(.A(n2585), .O(n2588));
  invx g2490(.A(n2555), .O(n2589));
  invx g2491(.A(n2559), .O(n2590));
  invx g2492(.A(n2744), .O(n2591));
  invx g2493(.A(n2744), .O(n2592));
  invx g2494(.A(n2584), .O(n2593));
  invx g2495(.A(n2564), .O(n2594));
  invx g2496(.A(n2542), .O(n2595));
  invx g2497(.A(n2579), .O(n2596));
  invx g2498(.A(n206), .O(n2597));
  invx g2499(.A(n202), .O(n2598));
  invx g2500(.A(n200), .O(n2599));
  invx g2501(.A(n198), .O(n2600));
  invx g2502(.A(n197), .O(n2601));
  invx g2503(.A(n196), .O(n2602));
  invx g2504(.A(n186), .O(n2603));
  invx g2505(.A(n185), .O(n2604));
  invx g2506(.A(n172), .O(n2605));
  invx g2507(.A(n163), .O(n2606));
  invx g2508(.A(n330), .O(n2607));
  invx g2509(.A(n1082), .O(n2608));
  invx g2510(.A(n1081), .O(n2609));
  invx g2511(.A(n584), .O(n2610));
  invx g2512(.A(n205), .O(n2611));
  invx g2513(.A(n1411), .O(n2612));
  invx g2514(.A(n299), .O(n2613));
  invx g2515(.A(n211), .O(n2614));
  invx g2516(.A(n294), .O(n2615));
  invx g2517(.A(n288), .O(n2616));
  invx g2518(.A(n329), .O(n2617));
  invx g2519(.A(n283), .O(n2618));
  invx g2520(.A(n284), .O(n2619));
  invx g2521(.A(n280), .O(n2620));
  invx g2522(.A(n276), .O(n2621));
  invx g2523(.A(n277), .O(n2622));
  invx g2524(.A(n683), .O(n2623));
  invx g2525(.A(n272), .O(n2624));
  invx g2526(.A(n266), .O(n2625));
  invx g2527(.A(n645), .O(n2626));
  invx g2528(.A(n711), .O(n2627));
  invx g2529(.A(n204), .O(n2628));
  invx g2530(.A(n267), .O(n2629));
  invx g2531(.A(n269), .O(n2630));
  invx g2532(.A(n261), .O(n2631));
  invx g2533(.A(n262), .O(n2632));
  invx g2534(.A(n1205), .O(n2633));
  invx g2535(.A(n248), .O(n2634));
  invx g2536(.A(n249), .O(n2635));
  invx g2537(.A(n244), .O(n2636));
  invx g2538(.A(n1162), .O(n2637));
  invx g2539(.A(n1161), .O(n2638));
  invx g2540(.A(n195), .O(n2639));
  invx g2541(.A(n210), .O(n2640));
  invx g2542(.A(n239), .O(n2641));
  invx g2543(.A(n233), .O(n2642));
  invx g2544(.A(n1136), .O(n2643));
  invx g2545(.A(n235), .O(n2644));
  invx g2546(.A(n236), .O(n2645));
  invx g2547(.A(n237), .O(n2646));
  invx g2548(.A(n224), .O(n2647));
  invx g2549(.A(n225), .O(n2648));
  invx g2550(.A(n228), .O(n2649));
  invx g2551(.A(n188), .O(n2650));
  invx g2552(.A(n229), .O(n2651));
  invx g2553(.A(n218), .O(n2652));
  invx g2554(.A(n217), .O(n2653));
  invx g2555(.A(n219), .O(n2654));
  invx g2556(.A(n221), .O(n2655));
  invx g2557(.A(n208), .O(n2656));
  invx g2558(.A(n212), .O(n2657));
  invx g2559(.A(n215), .O(n2658));
  invx g2560(.A(n214), .O(n2659));
  invx g2561(.A(n241), .O(n2660));
  invx g2562(.A(n553), .O(n2661));
  invx g2563(.A(n193), .O(n2662));
  invx g2564(.A(n187), .O(n2663));
  invx g2565(.A(n203), .O(n2664));
  invx g2566(.A(n201), .O(n2665));
  invx g2567(.A(n175), .O(n2666));
  invx g2568(.A(n199), .O(n2667));
  invx g2569(.A(n189), .O(n2668));
  invx g2570(.A(n856), .O(n2669));
  invx g2571(.A(n192), .O(n2670));
  invx g2572(.A(n190), .O(n2671));
  invx g2573(.A(n184), .O(n2672));
  invx g2574(.A(n176), .O(n2673));
  invx g2575(.A(n165), .O(n2674));
  invx g2576(.A(n182), .O(n2675));
  invx g2577(.A(n1928), .O(n2676));
  invx g2578(.A(n1518), .O(n2677));
  invx g2579(.A(n1533), .O(n2678));
  invx g2580(.A(n1513), .O(n2679));
  invx g2581(.A(n1516), .O(n2680));
  invx g2582(.A(n1506), .O(n2681));
  invx g2583(.A(n257), .O(n2682));
  invx g2584(.A(n2038), .O(n2683));
  invx g2585(.A(n776), .O(n2684));
  invx g2586(.A(n676), .O(n2685));
  invx g2587(.A(n1489), .O(n2686));
  invx g2588(.A(n1505), .O(n2687));
  invx g2589(.A(n2379), .O(n2688));
  invx g2590(.A(n2050), .O(n2689));
  invx g2591(.A(n1530), .O(n2690));
  invx g2592(.A(n1487), .O(n2691));
  invx g2593(.A(n1519), .O(n2692));
  invx g2594(.A(n1700), .O(n2693));
  invx g2595(.A(n650), .O(n2694));
  invx g2596(.A(n1541), .O(n2695));
  invx g2597(.A(n2048), .O(n2696));
  invx g2598(.A(n1566), .O(n2697));
  invx g2599(.A(n1507), .O(n2698));
  invx g2600(.A(n2386), .O(n2699));
  invx g2601(.A(n1554), .O(n2700));
  invx g2602(.A(n2049), .O(n2701));
  invx g2603(.A(n649), .O(n2702));
  invx g2604(.A(n1486), .O(n2703));
  invx g2605(.A(n1563), .O(n2704));
  invx g2606(.A(n1512), .O(n2705));
  invx g2607(.A(n1588), .O(n2706));
  invx g2608(.A(n1491), .O(n2707));
  invx g2609(.A(n1523), .O(n2708));
  invx g2610(.A(n2045), .O(n2709));
  invx g2611(.A(n2051), .O(n2710));
  invx g2612(.A(n596), .O(n2711));
  invx g2613(.A(n2046), .O(n2712));
  invx g2614(.A(n1550), .O(n2713));
  invx g2615(.A(n1540), .O(n2714));
  invx g2616(.A(n1503), .O(n2715));
  invx g2617(.A(n2076), .O(n2716));
  invx g2618(.A(n2078), .O(n2717));
  invx g2619(.A(n2392), .O(n2718));
  invx g2620(.A(n1643), .O(n2719));
  invx g2621(.A(n2058), .O(n2720));
  invx g2622(.A(n2053), .O(n2721));
  invx g2623(.A(n355), .O(n2722));
  invx g2624(.A(n1501), .O(n2723));
  invx g2625(.A(n1589), .O(n2724));
  invx g2626(.A(n1502), .O(n2725));
  invx g2627(.A(n1500), .O(n2726));
  invx g2628(.A(n1484), .O(n2727));
  invx g2629(.A(n1880), .O(n2728));
  invx g2630(.A(n328), .O(n2729));
  invx g2631(.A(n327), .O(n2730));
  invx g2632(.A(n354), .O(n2731));
  andx g2633(.A(n2733), .B(pi33), .O(n2732));
  andx g2634(.A(n2364), .B(n2734), .O(n2733));
  orx  g2635(.A(n2331), .B(n2735), .O(n2734));
  andx g2636(.A(n2736), .B(n2541), .O(n2735));
  orx  g2637(.A(n2738), .B(n2737), .O(n2736));
  orx  g2638(.A(n2454), .B(n2532), .O(n2737));
  andx g2639(.A(n2755), .B(n2361), .O(n2738));
  andx g2640(.A(n1587), .B(n2364), .O(n2739));
  andx g2641(.A(n1586), .B(n2402), .O(n2740));
  andx g2642(.A(n1585), .B(n2400), .O(n2741));
  andx g2643(.A(n2743), .B(n2375), .O(n2742));
  andx g2644(.A(n2745), .B(n2581), .O(n2743));
  invx g2645(.A(pi05), .O(n2744));
  orx  g2646(.A(n2761), .B(n2746), .O(n2745));
  andx g2647(.A(n2748), .B(n2351), .O(n2746));
  invx g2648(.A(pi06), .O(n2747));
  orx  g2649(.A(n2756), .B(n2749), .O(n2748));
  orx  g2650(.A(n2753), .B(n2750), .O(n2749));
  andx g2651(.A(n2752), .B(n2527), .O(n2750));
  invx g2652(.A(pi04), .O(n2751));
  invx g2653(.A(n2754), .O(n2752));
  andx g2654(.A(n2754), .B(pi04), .O(n2753));
  orx  g2655(.A(n2360), .B(n2755), .O(n2754));
  orx  g2656(.A(n2403), .B(n2357), .O(n2755));
  andx g2657(.A(n2758), .B(n2460), .O(n2756));
  invx g2658(.A(pi03), .O(n2757));
  orx  g2659(.A(n2759), .B(pi02), .O(n2758));
  andx g2660(.A(pi00), .B(n2356), .O(n2759));
  invx g2661(.A(pi01), .O(n2760));
  andx g2662(.A(n2766), .B(n2762), .O(n2761));
  andx g2663(.A(n2763), .B(pi03), .O(n2762));
  andx g2664(.A(n2440), .B(n2360), .O(n2763));
  invx g2665(.A(pi02), .O(n2764));
  invx g2666(.A(pi00), .O(n2765));
  andx g2667(.A(pi01), .B(pi04), .O(n2766));
  andx g2668(.A(n1584), .B(n2376), .O(n2767));
  andx g2669(.A(n1581), .B(n2367), .O(n2768));
  andx g2670(.A(n1578), .B(n2401), .O(n2769));
  andx g2671(.A(n1575), .B(n2374), .O(n2770));
  andx g2672(.A(n1573), .B(n2375), .O(n2771));
  andx g2673(.A(n1570), .B(n2819), .O(n2772));
  andx g2674(.A(n1568), .B(n2402), .O(n2773));
  andx g2675(.A(n1565), .B(n2400), .O(n2774));
  andx g2676(.A(n1562), .B(n2374), .O(n2775));
  andx g2677(.A(n1560), .B(n2376), .O(n2776));
  andx g2678(.A(n1558), .B(n2367), .O(n2777));
  andx g2679(.A(n1553), .B(n2401), .O(n2778));
  andx g2680(.A(n1549), .B(n2400), .O(n2779));
  andx g2681(.A(n1543), .B(n2375), .O(n2780));
  andx g2682(.A(n1539), .B(n2819), .O(n2781));
  andx g2683(.A(n1537), .B(n2402), .O(n2782));
  andx g2684(.A(n1532), .B(n2401), .O(n2783));
  andx g2685(.A(n1529), .B(n2374), .O(n2784));
  andx g2686(.A(n1526), .B(n2376), .O(n2785));
  andx g2687(.A(n1522), .B(n2367), .O(n2786));
  andx g2688(.A(n326), .B(n2402), .O(n2787));
  andx g2689(.A(n324), .B(n2400), .O(n2788));
  andx g2690(.A(n322), .B(n2375), .O(n2789));
  andx g2691(.A(n320), .B(n2364), .O(n2790));
  andx g2692(.A(n318), .B(n2364), .O(n2791));
  andx g2693(.A(n316), .B(n2401), .O(n2792));
  andx g2694(.A(n313), .B(n2374), .O(n2793));
  andx g2695(.A(n311), .B(n2376), .O(n2794));
  andx g2696(.A(n308), .B(n2364), .O(n2795));
  andx g2697(.A(n307), .B(n2402), .O(n2796));
  andx g2698(.A(n304), .B(n2400), .O(n2797));
  andx g2699(.A(n301), .B(n2375), .O(n2798));
  andx g2700(.A(n298), .B(n2376), .O(n2799));
  andx g2701(.A(n295), .B(n2367), .O(n2800));
  andx g2702(.A(n292), .B(n2401), .O(n2801));
  andx g2703(.A(n289), .B(n2374), .O(n2802));
  andx g2704(.A(n286), .B(n2375), .O(n2803));
  andx g2705(.A(n282), .B(n2364), .O(n2804));
  andx g2706(.A(n278), .B(n2402), .O(n2805));
  andx g2707(.A(n273), .B(n2400), .O(n2806));
  andx g2708(.A(n270), .B(n2374), .O(n2807));
  andx g2709(.A(n265), .B(n2376), .O(n2808));
  andx g2710(.A(n263), .B(n2367), .O(n2809));
  andx g2711(.A(n259), .B(n2401), .O(n2810));
  andx g2712(.A(n256), .B(n2400), .O(n2811));
  andx g2713(.A(n251), .B(n2375), .O(n2812));
  andx g2714(.A(n247), .B(n2819), .O(n2813));
  andx g2715(.A(n243), .B(n2402), .O(n2814));
  andx g2716(.A(n238), .B(n2401), .O(n2815));
  andx g2717(.A(n231), .B(n2374), .O(n2816));
  andx g2718(.A(n223), .B(n2376), .O(n2817));
  andx g2719(.A(n216), .B(n2367), .O(n2818));
  invx g2720(.A(n2820), .O(n2819));
  orx  g2721(.A(n2832), .B(n2821), .O(n2820));
  orx  g2722(.A(n2827), .B(n2822), .O(n2821));
  orx  g2723(.A(n2825), .B(n2823), .O(n2822));
  orx  g2724(.A(pi10), .B(n2824), .O(n2823));
  orx  g2725(.A(pi12), .B(pi11), .O(n2824));
  orx  g2726(.A(pi13), .B(n2826), .O(n2825));
  orx  g2727(.A(pi15), .B(pi14), .O(n2826));
  orx  g2728(.A(n2830), .B(n2828), .O(n2827));
  orx  g2729(.A(pi16), .B(n2829), .O(n2828));
  orx  g2730(.A(pi18), .B(pi17), .O(n2829));
  orx  g2731(.A(pi19), .B(n2831), .O(n2830));
  orx  g2732(.A(pi21), .B(pi20), .O(n2831));
  orx  g2733(.A(n2838), .B(n2833), .O(n2832));
  orx  g2734(.A(n2836), .B(n2834), .O(n2833));
  orx  g2735(.A(pi22), .B(n2835), .O(n2834));
  orx  g2736(.A(pi24), .B(pi23), .O(n2835));
  orx  g2737(.A(pi25), .B(n2837), .O(n2836));
  orx  g2738(.A(pi27), .B(pi26), .O(n2837));
  orx  g2739(.A(n2841), .B(n2839), .O(n2838));
  orx  g2740(.A(pi28), .B(n2840), .O(n2839));
  orx  g2741(.A(pi30), .B(pi29), .O(n2840));
  orx  g2742(.A(n2843), .B(n2842), .O(n2841));
  orx  g2743(.A(pi07), .B(pi31), .O(n2842));
  orx  g2744(.A(pi09), .B(pi08), .O(n2843));
endmodule


