// Benchmark "top" written by ABC on Fri Feb  7 13:49:46 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n172, n173, n174, n175, n176, n177, n178, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n191, n192, n194, n195,
    n196, n197, n198, n199, n200, n201, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n221,
    n222, n223, n224, n225, n226, n228, n229, n230, n231, n232, n233, n235,
    n236, n237, n238, n239, n240, n242, n243, n244, n245, n246, n247, n249,
    n250, n251, n252, n253, n254, n256, n257, n258, n259, n260, n261, n263,
    n264, n265, n266, n267, n268, n270, n271, n272, n273, n274, n275, n277,
    n278, n279, n280, n281, n282, n284, n285, n286, n287, n289, n290, n291,
    n292, n293, n294, n296, n297, n298, n299, n300, n301, n303, n304, n305,
    n306, n307, n308, n310, n311, n312, n313, n314, n315, n317, n318, n319,
    n320, n321, n322, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
    n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
    n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
    n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
    n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
    n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
    n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3491, n3492, n3493, n3494, n3495, n3496, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529;
  invx g0000(.A(n2930), .O(n64));
  invx g0001(.A(n64), .O(n65));
  invx g0002(.A(n2106), .O(n66));
  invx g0003(.A(n66), .O(n67));
  invx g0004(.A(n2640), .O(n68));
  invx g0005(.A(n68), .O(n69));
  invx g0006(.A(n138), .O(n70));
  invx g0007(.A(n70), .O(n71));
  invx g0008(.A(pi13), .O(n72));
  invx g0009(.A(pi11), .O(n73));
  invx g0010(.A(n1979), .O(n74));
  invx g0011(.A(n74), .O(n75));
  invx g0012(.A(n2298), .O(n76));
  invx g0013(.A(n76), .O(n77));
  invx g0014(.A(n2476), .O(n78));
  invx g0015(.A(n78), .O(n79));
  invx g0016(.A(n3049), .O(n80));
  invx g0017(.A(n80), .O(n81));
  invx g0018(.A(n3157), .O(n82));
  invx g0019(.A(n82), .O(n83));
  invx g0020(.A(n3255), .O(n84));
  invx g0021(.A(n84), .O(n85));
  invx g0022(.A(n3348), .O(n86));
  invx g0023(.A(n86), .O(n87));
  invx g0024(.A(n2790), .O(n88));
  invx g0025(.A(n88), .O(n89));
  invx g0026(.A(pi15), .O(n90));
  invx g0027(.A(pi01), .O(n91));
  invx g0028(.A(n3501), .O(n92));
  invx g0029(.A(n92), .O(n93));
  invx g0030(.A(pi13), .O(n94));
  invx g0031(.A(pi11), .O(n95));
  invx g0032(.A(pi11), .O(n96));
  invx g0033(.A(n1215), .O(n97));
  invx g0034(.A(n1215), .O(n98));
  invx g0035(.A(pi09), .O(n99));
  invx g0036(.A(pi09), .O(n100));
  invx g0037(.A(n1065), .O(n101));
  invx g0038(.A(n150), .O(n102));
  invx g0039(.A(pi07), .O(n103));
  invx g0040(.A(pi07), .O(n104));
  invx g0041(.A(pi05), .O(n105));
  invx g0042(.A(n138), .O(n106));
  invx g0043(.A(n106), .O(n107));
  invx g0044(.A(n106), .O(n108));
  invx g0045(.A(n184), .O(n109));
  invx g0046(.A(n185), .O(n110));
  invx g0047(.A(n183), .O(n111));
  invx g0048(.A(pi17), .O(n112));
  invx g0049(.A(pi17), .O(n113));
  invx g0050(.A(pi17), .O(n114));
  invx g0051(.A(pi17), .O(n115));
  invx g0052(.A(pi15), .O(n116));
  invx g0053(.A(pi15), .O(n117));
  invx g0054(.A(pi15), .O(n118));
  invx g0055(.A(pi15), .O(n119));
  invx g0056(.A(pi13), .O(n120));
  invx g0057(.A(pi13), .O(n121));
  invx g0058(.A(pi13), .O(n122));
  invx g0059(.A(pi01), .O(n123));
  invx g0060(.A(pi01), .O(n124));
  invx g0061(.A(pi01), .O(n125));
  invx g0062(.A(pi01), .O(n126));
  invx g0063(.A(pi11), .O(n127));
  invx g0064(.A(pi11), .O(n128));
  invx g0065(.A(pi11), .O(n129));
  invx g0066(.A(pi09), .O(n130));
  invx g0067(.A(pi09), .O(n131));
  invx g0068(.A(pi09), .O(n132));
  invx g0069(.A(pi07), .O(n133));
  invx g0070(.A(pi07), .O(n134));
  invx g0071(.A(pi07), .O(n135));
  invx g0072(.A(pi07), .O(n136));
  invx g0073(.A(pi05), .O(n137));
  invx g0074(.A(pi05), .O(n138));
  invx g0075(.A(pi05), .O(n139));
  bufx g0076(.A(n3529), .O(n140));
  bufx g0077(.A(n3528), .O(n141));
  bufx g0078(.A(n1584), .O(n142));
  bufx g0079(.A(n3527), .O(n143));
  bufx g0080(.A(n3527), .O(n144));
  invx g0081(.A(n97), .O(n145));
  invx g0082(.A(n98), .O(n146));
  bufx g0083(.A(n2764), .O(n147));
  bufx g0084(.A(n2612), .O(n148));
  bufx g0085(.A(n3139), .O(po16));
  bufx g0086(.A(n1065), .O(n150));
  bufx g0087(.A(n1065), .O(n151));
  bufx g0088(.A(n722), .O(n152));
  bufx g0089(.A(n722), .O(n153));
  bufx g0090(.A(n722), .O(n154));
  bufx g0091(.A(n1475), .O(n155));
  bufx g0092(.A(n1475), .O(n156));
  bufx g0093(.A(n2905), .O(n157));
  bufx g0094(.A(n2905), .O(n158));
  bufx g0095(.A(n2614), .O(n159));
  bufx g0096(.A(n2614), .O(po08));
  bufx g0097(.A(n2268), .O(po04));
  bufx g0098(.A(n2268), .O(n162));
  bufx g0099(.A(n2268), .O(n163));
  invx g0100(.A(pi03), .O(n164));
  bufx g0101(.A(n1759), .O(n165));
  bufx g0102(.A(n3236), .O(n166));
  bufx g0103(.A(n2446), .O(n167));
  bufx g0104(.A(n2446), .O(n168));
  bufx g0105(.A(n2072), .O(n169));
  bufx g0106(.A(n2072), .O(n170));
  bufx g0107(.A(n3029), .O(po14));
  bufx g0108(.A(n3029), .O(n172));
  bufx g0109(.A(n327), .O(n173));
  bufx g0110(.A(n327), .O(n174));
  bufx g0111(.A(n1353), .O(n175));
  bufx g0112(.A(n1353), .O(n176));
  bufx g0113(.A(n2266), .O(n177));
  bufx g0114(.A(n2266), .O(n178));
  bufx g0115(.A(n2766), .O(po10));
  bufx g0116(.A(n2766), .O(n180));
  bufx g0117(.A(n901), .O(n181));
  bufx g0118(.A(n901), .O(n182));
  bufx g0119(.A(n529), .O(n183));
  bufx g0120(.A(n529), .O(n184));
  bufx g0121(.A(n529), .O(n185));
  bufx g0122(.A(n1582), .O(n186));
  bufx g0123(.A(n3137), .O(n187));
  bufx g0124(.A(n1473), .O(n188));
  bufx g0125(.A(n3027), .O(n189));
  bufx g0126(.A(n3317), .O(po20));
  bufx g0127(.A(n1680), .O(n191));
  bufx g0128(.A(n1350), .O(n192));
  bufx g0129(.A(n2902), .O(po12));
  bufx g0130(.A(n899), .O(n194));
  bufx g0131(.A(n720), .O(n195));
  bufx g0132(.A(n720), .O(n196));
  bufx g0133(.A(n3526), .O(n197));
  bufx g0134(.A(n3526), .O(n198));
  bufx g0135(.A(n3526), .O(n199));
  bufx g0136(.A(po06), .O(n200));
  bufx g0137(.A(po06), .O(n201));
  bufx g0138(.A(n2074), .O(po02));
  bufx g0139(.A(n2074), .O(n203));
  bufx g0140(.A(n2074), .O(n204));
  bufx g0141(.A(n328), .O(n205));
  bufx g0142(.A(n328), .O(n206));
  bufx g0143(.A(n328), .O(n207));
  bufx g0144(.A(n3525), .O(n208));
  bufx g0145(.A(n3525), .O(n209));
  bufx g0146(.A(n3525), .O(n210));
  bufx g0147(.A(n3525), .O(n211));
  bufx g0148(.A(n3515), .O(n212));
  bufx g0149(.A(n3515), .O(n213));
  bufx g0150(.A(n3515), .O(n214));
  bufx g0151(.A(n3515), .O(n215));
  invx g0152(.A(pi03), .O(n216));
  invx g0153(.A(pi03), .O(n217));
  invx g0154(.A(pi03), .O(n218));
  invx g0155(.A(pi03), .O(n219));
  orx  g0156(.A(n222), .B(n221), .O(po19));
  andx g0157(.A(n173), .B(n455), .O(n221));
  andx g0158(.A(n223), .B(n206), .O(n222));
  orx  g0159(.A(n225), .B(n224), .O(n223));
  andx g0160(.A(n451), .B(n342), .O(n224));
  andx g0161(.A(n226), .B(n450), .O(n225));
  invx g0162(.A(n342), .O(n226));
  orx  g0163(.A(n229), .B(n228), .O(po17));
  andx g0164(.A(n174), .B(n443), .O(n228));
  andx g0165(.A(n230), .B(n207), .O(n229));
  orx  g0166(.A(n232), .B(n231), .O(n230));
  andx g0167(.A(n439), .B(n344), .O(n231));
  andx g0168(.A(n233), .B(n438), .O(n232));
  invx g0169(.A(n344), .O(n233));
  orx  g0170(.A(n236), .B(n235), .O(po15));
  andx g0171(.A(n327), .B(n431), .O(n235));
  andx g0172(.A(n237), .B(n207), .O(n236));
  orx  g0173(.A(n239), .B(n238), .O(n237));
  andx g0174(.A(n427), .B(n346), .O(n238));
  andx g0175(.A(n240), .B(n426), .O(n239));
  invx g0176(.A(n346), .O(n240));
  orx  g0177(.A(n243), .B(n242), .O(po13));
  andx g0178(.A(n173), .B(n419), .O(n242));
  andx g0179(.A(n244), .B(n206), .O(n243));
  orx  g0180(.A(n246), .B(n245), .O(n244));
  andx g0181(.A(n415), .B(n348), .O(n245));
  andx g0182(.A(n247), .B(n414), .O(n246));
  invx g0183(.A(n348), .O(n247));
  orx  g0184(.A(n250), .B(n249), .O(po11));
  andx g0185(.A(n174), .B(n407), .O(n249));
  andx g0186(.A(n251), .B(n207), .O(n250));
  orx  g0187(.A(n253), .B(n252), .O(n251));
  andx g0188(.A(n403), .B(n350), .O(n252));
  andx g0189(.A(n254), .B(n402), .O(n253));
  invx g0190(.A(n350), .O(n254));
  orx  g0191(.A(n257), .B(n256), .O(po09));
  andx g0192(.A(n174), .B(n395), .O(n256));
  andx g0193(.A(n258), .B(n205), .O(n257));
  orx  g0194(.A(n260), .B(n259), .O(n258));
  andx g0195(.A(n391), .B(n352), .O(n259));
  andx g0196(.A(n261), .B(n390), .O(n260));
  invx g0197(.A(n352), .O(n261));
  orx  g0198(.A(n264), .B(n263), .O(po07));
  andx g0199(.A(n173), .B(n383), .O(n263));
  andx g0200(.A(n265), .B(n206), .O(n264));
  orx  g0201(.A(n267), .B(n266), .O(n265));
  andx g0202(.A(n379), .B(n354), .O(n266));
  andx g0203(.A(n268), .B(n378), .O(n267));
  invx g0204(.A(n354), .O(n268));
  orx  g0205(.A(n271), .B(n270), .O(po05));
  andx g0206(.A(n174), .B(n372), .O(n270));
  andx g0207(.A(n272), .B(n207), .O(n271));
  orx  g0208(.A(n274), .B(n273), .O(n272));
  andx g0209(.A(n368), .B(n356), .O(n273));
  andx g0210(.A(n275), .B(n367), .O(n274));
  invx g0211(.A(n356), .O(n275));
  orx  g0212(.A(n282), .B(n277), .O(po03));
  andx g0213(.A(n278), .B(n207), .O(n277));
  andx g0214(.A(n280), .B(n279), .O(n278));
  orx  g0215(.A(n75), .B(n359), .O(n279));
  orx  g0216(.A(n74), .B(n281), .O(n280));
  invx g0217(.A(n359), .O(n281));
  andx g0218(.A(n327), .B(n363), .O(n282));
  orx  g0219(.A(n285), .B(n284), .O(po31));
  andx g0220(.A(n173), .B(n526), .O(n284));
  andx g0221(.A(n286), .B(n206), .O(n285));
  andx g0222(.A(n287), .B(n330), .O(n286));
  invx g0223(.A(n522), .O(n287));
  orx  g0224(.A(n290), .B(n289), .O(po29));
  andx g0225(.A(n174), .B(n515), .O(n289));
  andx g0226(.A(n291), .B(n207), .O(n290));
  orx  g0227(.A(n293), .B(n292), .O(n291));
  andx g0228(.A(n511), .B(n332), .O(n292));
  andx g0229(.A(n294), .B(n510), .O(n293));
  invx g0230(.A(n332), .O(n294));
  orx  g0231(.A(n297), .B(n296), .O(po27));
  andx g0232(.A(n327), .B(n503), .O(n296));
  andx g0233(.A(n298), .B(n328), .O(n297));
  orx  g0234(.A(n300), .B(n299), .O(n298));
  andx g0235(.A(n499), .B(n334), .O(n299));
  andx g0236(.A(n301), .B(n498), .O(n300));
  invx g0237(.A(n334), .O(n301));
  orx  g0238(.A(n304), .B(n303), .O(po25));
  andx g0239(.A(n173), .B(n491), .O(n303));
  andx g0240(.A(n305), .B(n206), .O(n304));
  orx  g0241(.A(n307), .B(n306), .O(n305));
  andx g0242(.A(n487), .B(n336), .O(n306));
  andx g0243(.A(n308), .B(n486), .O(n307));
  invx g0244(.A(n336), .O(n308));
  orx  g0245(.A(n311), .B(n310), .O(po23));
  andx g0246(.A(n174), .B(n479), .O(n310));
  andx g0247(.A(n312), .B(n205), .O(n311));
  orx  g0248(.A(n314), .B(n313), .O(n312));
  andx g0249(.A(n475), .B(n338), .O(n313));
  andx g0250(.A(n315), .B(n474), .O(n314));
  invx g0251(.A(n338), .O(n315));
  orx  g0252(.A(n318), .B(n317), .O(po21));
  andx g0253(.A(n327), .B(n467), .O(n317));
  andx g0254(.A(n319), .B(n205), .O(n318));
  orx  g0255(.A(n321), .B(n320), .O(n319));
  andx g0256(.A(n463), .B(n340), .O(n320));
  andx g0257(.A(n322), .B(n462), .O(n321));
  invx g0258(.A(n340), .O(n322));
  orx  g0259(.A(n325), .B(n324), .O(po01));
  andx g0260(.A(n74), .B(n205), .O(n324));
  andx g0261(.A(pi00), .B(n326), .O(n325));
  orx  g0262(.A(n173), .B(n123), .O(n326));
  invx g0263(.A(n205), .O(n327));
  orx  g0264(.A(n329), .B(n524), .O(n328));
  andx g0265(.A(n522), .B(n330), .O(n329));
  orx  g0266(.A(n331), .B(n512), .O(n330));
  andx g0267(.A(n510), .B(n332), .O(n331));
  orx  g0268(.A(n333), .B(n500), .O(n332));
  andx g0269(.A(n498), .B(n334), .O(n333));
  orx  g0270(.A(n335), .B(n488), .O(n334));
  andx g0271(.A(n486), .B(n336), .O(n335));
  orx  g0272(.A(n337), .B(n476), .O(n336));
  andx g0273(.A(n474), .B(n338), .O(n337));
  orx  g0274(.A(n339), .B(n464), .O(n338));
  andx g0275(.A(n462), .B(n340), .O(n339));
  orx  g0276(.A(n341), .B(n452), .O(n340));
  andx g0277(.A(n450), .B(n342), .O(n341));
  orx  g0278(.A(n343), .B(n440), .O(n342));
  andx g0279(.A(n438), .B(n344), .O(n343));
  orx  g0280(.A(n345), .B(n428), .O(n344));
  andx g0281(.A(n426), .B(n346), .O(n345));
  orx  g0282(.A(n347), .B(n416), .O(n346));
  andx g0283(.A(n414), .B(n348), .O(n347));
  orx  g0284(.A(n349), .B(n404), .O(n348));
  andx g0285(.A(n402), .B(n350), .O(n349));
  orx  g0286(.A(n351), .B(n392), .O(n350));
  andx g0287(.A(n390), .B(n352), .O(n351));
  orx  g0288(.A(n353), .B(n380), .O(n352));
  andx g0289(.A(n378), .B(n354), .O(n353));
  orx  g0290(.A(n355), .B(n369), .O(n354));
  andx g0291(.A(n367), .B(n356), .O(n355));
  orx  g0292(.A(n358), .B(n357), .O(n356));
  andx g0293(.A(n363), .B(n216), .O(n357));
  andx g0294(.A(n359), .B(n75), .O(n358));
  orx  g0295(.A(n362), .B(n360), .O(n359));
  invx g0296(.A(n361), .O(n360));
  orx  g0297(.A(n363), .B(pi03), .O(n361));
  andx g0298(.A(pi03), .B(n363), .O(n362));
  orx  g0299(.A(n365), .B(n364), .O(n363));
  andx g0300(.A(n66), .B(n185), .O(n364));
  andx g0301(.A(pi02), .B(n366), .O(n365));
  orx  g0302(.A(n109), .B(n91), .O(n366));
  invx g0303(.A(n368), .O(n367));
  orx  g0304(.A(n370), .B(n369), .O(n368));
  andx g0305(.A(n372), .B(n3518), .O(n369));
  invx g0306(.A(n371), .O(n370));
  orx  g0307(.A(n372), .B(n105), .O(n371));
  orx  g0308(.A(n377), .B(n373), .O(n372));
  andx g0309(.A(n374), .B(n184), .O(n373));
  andx g0310(.A(n376), .B(n375), .O(n374));
  orx  g0311(.A(n67), .B(n561), .O(n375));
  orx  g0312(.A(n66), .B(n562), .O(n376));
  andx g0313(.A(n111), .B(n566), .O(n377));
  invx g0314(.A(n379), .O(n378));
  orx  g0315(.A(n381), .B(n380), .O(n379));
  andx g0316(.A(n383), .B(n136), .O(n380));
  invx g0317(.A(n382), .O(n381));
  orx  g0318(.A(n383), .B(n133), .O(n382));
  orx  g0319(.A(n385), .B(n384), .O(n383));
  andx g0320(.A(n110), .B(n575), .O(n384));
  andx g0321(.A(n386), .B(n184), .O(n385));
  orx  g0322(.A(n388), .B(n387), .O(n386));
  andx g0323(.A(n571), .B(n558), .O(n387));
  andx g0324(.A(n389), .B(n570), .O(n388));
  invx g0325(.A(n558), .O(n389));
  invx g0326(.A(n391), .O(n390));
  orx  g0327(.A(n393), .B(n392), .O(n391));
  andx g0328(.A(n395), .B(n3522), .O(n392));
  invx g0329(.A(n394), .O(n393));
  orx  g0330(.A(n395), .B(n3522), .O(n394));
  orx  g0331(.A(n397), .B(n396), .O(n395));
  andx g0332(.A(n109), .B(n586), .O(n396));
  andx g0333(.A(n398), .B(n183), .O(n397));
  orx  g0334(.A(n400), .B(n399), .O(n398));
  andx g0335(.A(n582), .B(n556), .O(n399));
  andx g0336(.A(n401), .B(n581), .O(n400));
  invx g0337(.A(n556), .O(n401));
  invx g0338(.A(n403), .O(n402));
  orx  g0339(.A(n405), .B(n404), .O(n403));
  andx g0340(.A(n407), .B(n96), .O(n404));
  invx g0341(.A(n406), .O(n405));
  orx  g0342(.A(n95), .B(n407), .O(n406));
  orx  g0343(.A(n409), .B(n408), .O(n407));
  andx g0344(.A(n111), .B(n598), .O(n408));
  andx g0345(.A(n410), .B(n185), .O(n409));
  orx  g0346(.A(n412), .B(n411), .O(n410));
  andx g0347(.A(n594), .B(n554), .O(n411));
  andx g0348(.A(n413), .B(n593), .O(n412));
  invx g0349(.A(n554), .O(n413));
  invx g0350(.A(n415), .O(n414));
  orx  g0351(.A(n417), .B(n416), .O(n415));
  andx g0352(.A(n419), .B(n72), .O(n416));
  invx g0353(.A(n418), .O(n417));
  orx  g0354(.A(n121), .B(n419), .O(n418));
  orx  g0355(.A(n421), .B(n420), .O(n419));
  andx g0356(.A(n110), .B(n610), .O(n420));
  andx g0357(.A(n422), .B(n184), .O(n421));
  orx  g0358(.A(n424), .B(n423), .O(n422));
  andx g0359(.A(n606), .B(n552), .O(n423));
  andx g0360(.A(n425), .B(n605), .O(n424));
  invx g0361(.A(n552), .O(n425));
  invx g0362(.A(n427), .O(n426));
  orx  g0363(.A(n429), .B(n428), .O(n427));
  andx g0364(.A(n431), .B(n119), .O(n428));
  invx g0365(.A(n430), .O(n429));
  orx  g0366(.A(n90), .B(n431), .O(n430));
  orx  g0367(.A(n433), .B(n432), .O(n431));
  andx g0368(.A(n109), .B(n622), .O(n432));
  andx g0369(.A(n434), .B(n185), .O(n433));
  orx  g0370(.A(n436), .B(n435), .O(n434));
  andx g0371(.A(n618), .B(n550), .O(n435));
  andx g0372(.A(n437), .B(n617), .O(n436));
  invx g0373(.A(n550), .O(n437));
  invx g0374(.A(n439), .O(n438));
  orx  g0375(.A(n441), .B(n440), .O(n439));
  andx g0376(.A(n443), .B(n115), .O(n440));
  invx g0377(.A(n442), .O(n441));
  orx  g0378(.A(n3524), .B(n443), .O(n442));
  orx  g0379(.A(n445), .B(n444), .O(n443));
  andx g0380(.A(n111), .B(n634), .O(n444));
  andx g0381(.A(n446), .B(n183), .O(n445));
  orx  g0382(.A(n448), .B(n447), .O(n446));
  andx g0383(.A(n630), .B(n548), .O(n447));
  andx g0384(.A(n449), .B(n629), .O(n448));
  invx g0385(.A(n548), .O(n449));
  invx g0386(.A(n451), .O(n450));
  orx  g0387(.A(n453), .B(n452), .O(n451));
  andx g0388(.A(n455), .B(n212), .O(n452));
  invx g0389(.A(n454), .O(n453));
  orx  g0390(.A(n214), .B(n455), .O(n454));
  orx  g0391(.A(n457), .B(n456), .O(n455));
  andx g0392(.A(n110), .B(n646), .O(n456));
  andx g0393(.A(n458), .B(n185), .O(n457));
  orx  g0394(.A(n460), .B(n459), .O(n458));
  andx g0395(.A(n642), .B(n546), .O(n459));
  andx g0396(.A(n461), .B(n641), .O(n460));
  invx g0397(.A(n546), .O(n461));
  invx g0398(.A(n463), .O(n462));
  orx  g0399(.A(n465), .B(n464), .O(n463));
  andx g0400(.A(n467), .B(n210), .O(n464));
  invx g0401(.A(n466), .O(n465));
  orx  g0402(.A(n210), .B(n467), .O(n466));
  orx  g0403(.A(n469), .B(n468), .O(n467));
  andx g0404(.A(n109), .B(n658), .O(n468));
  andx g0405(.A(n470), .B(n184), .O(n469));
  orx  g0406(.A(n472), .B(n471), .O(n470));
  andx g0407(.A(n654), .B(n544), .O(n471));
  andx g0408(.A(n473), .B(n653), .O(n472));
  invx g0409(.A(n544), .O(n473));
  invx g0410(.A(n475), .O(n474));
  orx  g0411(.A(n477), .B(n476), .O(n475));
  andx g0412(.A(n479), .B(n197), .O(n476));
  invx g0413(.A(n478), .O(n477));
  orx  g0414(.A(n199), .B(n479), .O(n478));
  orx  g0415(.A(n481), .B(n480), .O(n479));
  andx g0416(.A(n111), .B(n670), .O(n480));
  andx g0417(.A(n482), .B(n183), .O(n481));
  orx  g0418(.A(n484), .B(n483), .O(n482));
  andx g0419(.A(n666), .B(n542), .O(n483));
  andx g0420(.A(n485), .B(n665), .O(n484));
  invx g0421(.A(n542), .O(n485));
  invx g0422(.A(n487), .O(n486));
  orx  g0423(.A(n489), .B(n488), .O(n487));
  andx g0424(.A(n491), .B(n144), .O(n488));
  invx g0425(.A(n490), .O(n489));
  orx  g0426(.A(n143), .B(n491), .O(n490));
  orx  g0427(.A(n493), .B(n492), .O(n491));
  andx g0428(.A(n110), .B(n682), .O(n492));
  andx g0429(.A(n494), .B(n183), .O(n493));
  orx  g0430(.A(n496), .B(n495), .O(n494));
  andx g0431(.A(n678), .B(n540), .O(n495));
  andx g0432(.A(n497), .B(n677), .O(n496));
  invx g0433(.A(n540), .O(n497));
  invx g0434(.A(n499), .O(n498));
  orx  g0435(.A(n501), .B(n500), .O(n499));
  andx g0436(.A(n503), .B(n141), .O(n500));
  invx g0437(.A(n502), .O(n501));
  orx  g0438(.A(n3528), .B(n503), .O(n502));
  orx  g0439(.A(n505), .B(n504), .O(n503));
  andx g0440(.A(n109), .B(n694), .O(n504));
  andx g0441(.A(n506), .B(n185), .O(n505));
  orx  g0442(.A(n508), .B(n507), .O(n506));
  andx g0443(.A(n690), .B(n538), .O(n507));
  andx g0444(.A(n509), .B(n689), .O(n508));
  invx g0445(.A(n538), .O(n509));
  invx g0446(.A(n511), .O(n510));
  orx  g0447(.A(n513), .B(n512), .O(n511));
  andx g0448(.A(n515), .B(n140), .O(n512));
  invx g0449(.A(n514), .O(n513));
  orx  g0450(.A(n3529), .B(n515), .O(n514));
  orx  g0451(.A(n517), .B(n516), .O(n515));
  andx g0452(.A(n111), .B(n706), .O(n516));
  andx g0453(.A(n518), .B(n184), .O(n517));
  orx  g0454(.A(n520), .B(n519), .O(n518));
  andx g0455(.A(n702), .B(n536), .O(n519));
  andx g0456(.A(n521), .B(n701), .O(n520));
  invx g0457(.A(n536), .O(n521));
  andx g0458(.A(n525), .B(n523), .O(n522));
  invx g0459(.A(n524), .O(n523));
  andx g0460(.A(n526), .B(n3514), .O(n524));
  orx  g0461(.A(n3514), .B(n526), .O(n525));
  orx  g0462(.A(n528), .B(n527), .O(n526));
  andx g0463(.A(n110), .B(n718), .O(n527));
  andx g0464(.A(n533), .B(n529), .O(n528));
  orx  g0465(.A(n531), .B(n530), .O(n529));
  andx g0466(.A(n3513), .B(n718), .O(n530));
  andx g0467(.A(n532), .B(n714), .O(n531));
  andx g0468(.A(n534), .B(n3514), .O(n532));
  andx g0469(.A(n713), .B(n534), .O(n533));
  orx  g0470(.A(n535), .B(n703), .O(n534));
  andx g0471(.A(n701), .B(n536), .O(n535));
  orx  g0472(.A(n537), .B(n691), .O(n536));
  andx g0473(.A(n689), .B(n538), .O(n537));
  orx  g0474(.A(n539), .B(n679), .O(n538));
  andx g0475(.A(n677), .B(n540), .O(n539));
  orx  g0476(.A(n541), .B(n667), .O(n540));
  andx g0477(.A(n665), .B(n542), .O(n541));
  orx  g0478(.A(n543), .B(n655), .O(n542));
  andx g0479(.A(n653), .B(n544), .O(n543));
  orx  g0480(.A(n545), .B(n643), .O(n544));
  andx g0481(.A(n641), .B(n546), .O(n545));
  orx  g0482(.A(n547), .B(n631), .O(n546));
  andx g0483(.A(n629), .B(n548), .O(n547));
  orx  g0484(.A(n549), .B(n619), .O(n548));
  andx g0485(.A(n617), .B(n550), .O(n549));
  orx  g0486(.A(n551), .B(n607), .O(n550));
  andx g0487(.A(n605), .B(n552), .O(n551));
  orx  g0488(.A(n553), .B(n595), .O(n552));
  andx g0489(.A(n593), .B(n554), .O(n553));
  orx  g0490(.A(n555), .B(n583), .O(n554));
  andx g0491(.A(n581), .B(n556), .O(n555));
  orx  g0492(.A(n557), .B(n572), .O(n556));
  andx g0493(.A(n570), .B(n558), .O(n557));
  orx  g0494(.A(n560), .B(n559), .O(n558));
  andx g0495(.A(n566), .B(n164), .O(n559));
  andx g0496(.A(n561), .B(n67), .O(n560));
  invx g0497(.A(n562), .O(n561));
  andx g0498(.A(n564), .B(n563), .O(n562));
  orx  g0499(.A(n566), .B(pi03), .O(n563));
  invx g0500(.A(n565), .O(n564));
  andx g0501(.A(pi03), .B(n566), .O(n565));
  orx  g0502(.A(n568), .B(n567), .O(n566));
  andx g0503(.A(n76), .B(n154), .O(n567));
  andx g0504(.A(pi04), .B(n569), .O(n568));
  orx  g0505(.A(n195), .B(n124), .O(n569));
  invx g0506(.A(n571), .O(n570));
  orx  g0507(.A(n573), .B(n572), .O(n571));
  andx g0508(.A(n107), .B(n575), .O(n572));
  invx g0509(.A(n574), .O(n573));
  orx  g0510(.A(n575), .B(n107), .O(n574));
  orx  g0511(.A(n580), .B(n576), .O(n575));
  andx g0512(.A(n577), .B(n153), .O(n576));
  andx g0513(.A(n579), .B(n578), .O(n577));
  orx  g0514(.A(n77), .B(n752), .O(n578));
  orx  g0515(.A(n76), .B(n753), .O(n579));
  andx g0516(.A(n196), .B(n757), .O(n580));
  invx g0517(.A(n582), .O(n581));
  orx  g0518(.A(n584), .B(n583), .O(n582));
  andx g0519(.A(n586), .B(n104), .O(n583));
  invx g0520(.A(n585), .O(n584));
  orx  g0521(.A(n586), .B(n104), .O(n585));
  orx  g0522(.A(n588), .B(n587), .O(n586));
  andx g0523(.A(n195), .B(n766), .O(n587));
  andx g0524(.A(n589), .B(n152), .O(n588));
  orx  g0525(.A(n591), .B(n590), .O(n589));
  andx g0526(.A(n762), .B(n749), .O(n590));
  andx g0527(.A(n592), .B(n761), .O(n591));
  invx g0528(.A(n749), .O(n592));
  invx g0529(.A(n594), .O(n593));
  orx  g0530(.A(n596), .B(n595), .O(n594));
  andx g0531(.A(n598), .B(n132), .O(n595));
  invx g0532(.A(n597), .O(n596));
  orx  g0533(.A(n598), .B(n131), .O(n597));
  orx  g0534(.A(n600), .B(n599), .O(n598));
  andx g0535(.A(n196), .B(n777), .O(n599));
  andx g0536(.A(n601), .B(n154), .O(n600));
  orx  g0537(.A(n603), .B(n602), .O(n601));
  andx g0538(.A(n773), .B(n747), .O(n602));
  andx g0539(.A(n604), .B(n772), .O(n603));
  invx g0540(.A(n747), .O(n604));
  invx g0541(.A(n606), .O(n605));
  orx  g0542(.A(n608), .B(n607), .O(n606));
  andx g0543(.A(n610), .B(n129), .O(n607));
  invx g0544(.A(n609), .O(n608));
  orx  g0545(.A(n73), .B(n610), .O(n609));
  orx  g0546(.A(n612), .B(n611), .O(n610));
  andx g0547(.A(n195), .B(n789), .O(n611));
  andx g0548(.A(n613), .B(n153), .O(n612));
  orx  g0549(.A(n615), .B(n614), .O(n613));
  andx g0550(.A(n785), .B(n745), .O(n614));
  andx g0551(.A(n616), .B(n784), .O(n615));
  invx g0552(.A(n745), .O(n616));
  invx g0553(.A(n618), .O(n617));
  orx  g0554(.A(n620), .B(n619), .O(n618));
  andx g0555(.A(n622), .B(n120), .O(n619));
  invx g0556(.A(n621), .O(n620));
  orx  g0557(.A(n94), .B(n622), .O(n621));
  orx  g0558(.A(n624), .B(n623), .O(n622));
  andx g0559(.A(n196), .B(n801), .O(n623));
  andx g0560(.A(n625), .B(n152), .O(n624));
  orx  g0561(.A(n627), .B(n626), .O(n625));
  andx g0562(.A(n797), .B(n743), .O(n626));
  andx g0563(.A(n628), .B(n796), .O(n627));
  invx g0564(.A(n743), .O(n628));
  invx g0565(.A(n630), .O(n629));
  orx  g0566(.A(n632), .B(n631), .O(n630));
  andx g0567(.A(n634), .B(n117), .O(n631));
  invx g0568(.A(n633), .O(n632));
  orx  g0569(.A(n118), .B(n634), .O(n633));
  orx  g0570(.A(n636), .B(n635), .O(n634));
  andx g0571(.A(n195), .B(n813), .O(n635));
  andx g0572(.A(n637), .B(n154), .O(n636));
  orx  g0573(.A(n639), .B(n638), .O(n637));
  andx g0574(.A(n809), .B(n741), .O(n638));
  andx g0575(.A(n640), .B(n808), .O(n639));
  invx g0576(.A(n741), .O(n640));
  invx g0577(.A(n642), .O(n641));
  orx  g0578(.A(n644), .B(n643), .O(n642));
  andx g0579(.A(n646), .B(n112), .O(n643));
  invx g0580(.A(n645), .O(n644));
  orx  g0581(.A(n113), .B(n646), .O(n645));
  orx  g0582(.A(n648), .B(n647), .O(n646));
  andx g0583(.A(n196), .B(n825), .O(n647));
  andx g0584(.A(n649), .B(n153), .O(n648));
  orx  g0585(.A(n651), .B(n650), .O(n649));
  andx g0586(.A(n821), .B(n739), .O(n650));
  andx g0587(.A(n652), .B(n820), .O(n651));
  invx g0588(.A(n739), .O(n652));
  invx g0589(.A(n654), .O(n653));
  orx  g0590(.A(n656), .B(n655), .O(n654));
  andx g0591(.A(n658), .B(n215), .O(n655));
  invx g0592(.A(n657), .O(n656));
  orx  g0593(.A(n213), .B(n658), .O(n657));
  orx  g0594(.A(n660), .B(n659), .O(n658));
  andx g0595(.A(n195), .B(n837), .O(n659));
  andx g0596(.A(n661), .B(n152), .O(n660));
  orx  g0597(.A(n663), .B(n662), .O(n661));
  andx g0598(.A(n833), .B(n737), .O(n662));
  andx g0599(.A(n664), .B(n832), .O(n663));
  invx g0600(.A(n737), .O(n664));
  invx g0601(.A(n666), .O(n665));
  orx  g0602(.A(n668), .B(n667), .O(n666));
  andx g0603(.A(n670), .B(n209), .O(n667));
  invx g0604(.A(n669), .O(n668));
  orx  g0605(.A(n209), .B(n670), .O(n669));
  orx  g0606(.A(n672), .B(n671), .O(n670));
  andx g0607(.A(n196), .B(n849), .O(n671));
  andx g0608(.A(n673), .B(n154), .O(n672));
  orx  g0609(.A(n675), .B(n674), .O(n673));
  andx g0610(.A(n845), .B(n735), .O(n674));
  andx g0611(.A(n676), .B(n844), .O(n675));
  invx g0612(.A(n735), .O(n676));
  invx g0613(.A(n678), .O(n677));
  orx  g0614(.A(n680), .B(n679), .O(n678));
  andx g0615(.A(n682), .B(n199), .O(n679));
  invx g0616(.A(n681), .O(n680));
  orx  g0617(.A(n198), .B(n682), .O(n681));
  orx  g0618(.A(n684), .B(n683), .O(n682));
  andx g0619(.A(n195), .B(n861), .O(n683));
  andx g0620(.A(n685), .B(n153), .O(n684));
  orx  g0621(.A(n687), .B(n686), .O(n685));
  andx g0622(.A(n857), .B(n733), .O(n686));
  andx g0623(.A(n688), .B(n856), .O(n687));
  invx g0624(.A(n733), .O(n688));
  invx g0625(.A(n690), .O(n689));
  orx  g0626(.A(n692), .B(n691), .O(n690));
  andx g0627(.A(n694), .B(n3527), .O(n691));
  invx g0628(.A(n693), .O(n692));
  orx  g0629(.A(n144), .B(n694), .O(n693));
  orx  g0630(.A(n696), .B(n695), .O(n694));
  andx g0631(.A(n196), .B(n873), .O(n695));
  andx g0632(.A(n697), .B(n152), .O(n696));
  orx  g0633(.A(n699), .B(n698), .O(n697));
  andx g0634(.A(n869), .B(n731), .O(n698));
  andx g0635(.A(n700), .B(n868), .O(n699));
  invx g0636(.A(n731), .O(n700));
  invx g0637(.A(n702), .O(n701));
  orx  g0638(.A(n704), .B(n703), .O(n702));
  andx g0639(.A(n706), .B(n141), .O(n703));
  invx g0640(.A(n705), .O(n704));
  orx  g0641(.A(n3528), .B(n706), .O(n705));
  orx  g0642(.A(n708), .B(n707), .O(n706));
  andx g0643(.A(n195), .B(n885), .O(n707));
  andx g0644(.A(n709), .B(n154), .O(n708));
  orx  g0645(.A(n711), .B(n710), .O(n709));
  andx g0646(.A(n881), .B(n729), .O(n710));
  andx g0647(.A(n712), .B(n880), .O(n711));
  invx g0648(.A(n729), .O(n712));
  invx g0649(.A(n714), .O(n713));
  andx g0650(.A(n717), .B(n715), .O(n714));
  invx g0651(.A(n716), .O(n715));
  andx g0652(.A(n718), .B(n140), .O(n716));
  orx  g0653(.A(n3529), .B(n718), .O(n717));
  orx  g0654(.A(n721), .B(n719), .O(n718));
  andx g0655(.A(n196), .B(n897), .O(n719));
  invx g0656(.A(n152), .O(n720));
  andx g0657(.A(n726), .B(n153), .O(n721));
  orx  g0658(.A(n724), .B(n723), .O(n722));
  andx g0659(.A(n3512), .B(n897), .O(n723));
  andx g0660(.A(n725), .B(n893), .O(n724));
  andx g0661(.A(n3513), .B(n727), .O(n725));
  andx g0662(.A(n892), .B(n727), .O(n726));
  orx  g0663(.A(n728), .B(n882), .O(n727));
  andx g0664(.A(n880), .B(n729), .O(n728));
  orx  g0665(.A(n730), .B(n870), .O(n729));
  andx g0666(.A(n868), .B(n731), .O(n730));
  orx  g0667(.A(n732), .B(n858), .O(n731));
  andx g0668(.A(n856), .B(n733), .O(n732));
  orx  g0669(.A(n734), .B(n846), .O(n733));
  andx g0670(.A(n844), .B(n735), .O(n734));
  orx  g0671(.A(n736), .B(n834), .O(n735));
  andx g0672(.A(n832), .B(n737), .O(n736));
  orx  g0673(.A(n738), .B(n822), .O(n737));
  andx g0674(.A(n820), .B(n739), .O(n738));
  orx  g0675(.A(n740), .B(n810), .O(n739));
  andx g0676(.A(n808), .B(n741), .O(n740));
  orx  g0677(.A(n742), .B(n798), .O(n741));
  andx g0678(.A(n796), .B(n743), .O(n742));
  orx  g0679(.A(n744), .B(n786), .O(n743));
  andx g0680(.A(n784), .B(n745), .O(n744));
  orx  g0681(.A(n746), .B(n774), .O(n745));
  andx g0682(.A(n772), .B(n747), .O(n746));
  orx  g0683(.A(n748), .B(n763), .O(n747));
  andx g0684(.A(n761), .B(n749), .O(n748));
  orx  g0685(.A(n751), .B(n750), .O(n749));
  andx g0686(.A(n757), .B(n219), .O(n750));
  andx g0687(.A(n752), .B(n77), .O(n751));
  invx g0688(.A(n753), .O(n752));
  andx g0689(.A(n755), .B(n754), .O(n753));
  orx  g0690(.A(n757), .B(pi03), .O(n754));
  invx g0691(.A(n756), .O(n755));
  andx g0692(.A(pi03), .B(n757), .O(n756));
  orx  g0693(.A(n759), .B(n758), .O(n757));
  andx g0694(.A(n78), .B(n182), .O(n758));
  andx g0695(.A(pi06), .B(n760), .O(n759));
  orx  g0696(.A(n899), .B(n124), .O(n760));
  invx g0697(.A(n762), .O(n761));
  orx  g0698(.A(n764), .B(n763), .O(n762));
  andx g0699(.A(n766), .B(n3518), .O(n763));
  invx g0700(.A(n765), .O(n764));
  orx  g0701(.A(n766), .B(n137), .O(n765));
  orx  g0702(.A(n771), .B(n767), .O(n766));
  andx g0703(.A(n768), .B(n181), .O(n767));
  andx g0704(.A(n770), .B(n769), .O(n768));
  orx  g0705(.A(n79), .B(n929), .O(n769));
  orx  g0706(.A(n78), .B(n930), .O(n770));
  andx g0707(.A(n899), .B(n934), .O(n771));
  invx g0708(.A(n773), .O(n772));
  orx  g0709(.A(n775), .B(n774), .O(n773));
  andx g0710(.A(n777), .B(n136), .O(n774));
  invx g0711(.A(n776), .O(n775));
  orx  g0712(.A(n777), .B(n136), .O(n776));
  orx  g0713(.A(n779), .B(n778), .O(n777));
  andx g0714(.A(n194), .B(n943), .O(n778));
  andx g0715(.A(n780), .B(n182), .O(n779));
  orx  g0716(.A(n782), .B(n781), .O(n780));
  andx g0717(.A(n939), .B(n926), .O(n781));
  andx g0718(.A(n783), .B(n938), .O(n782));
  invx g0719(.A(n926), .O(n783));
  invx g0720(.A(n785), .O(n784));
  orx  g0721(.A(n787), .B(n786), .O(n785));
  andx g0722(.A(n789), .B(n3522), .O(n786));
  invx g0723(.A(n788), .O(n787));
  orx  g0724(.A(n789), .B(n99), .O(n788));
  orx  g0725(.A(n791), .B(n790), .O(n789));
  andx g0726(.A(n194), .B(n954), .O(n790));
  andx g0727(.A(n792), .B(n181), .O(n791));
  orx  g0728(.A(n794), .B(n793), .O(n792));
  andx g0729(.A(n950), .B(n924), .O(n793));
  andx g0730(.A(n795), .B(n949), .O(n794));
  invx g0731(.A(n924), .O(n795));
  invx g0732(.A(n797), .O(n796));
  orx  g0733(.A(n799), .B(n798), .O(n797));
  andx g0734(.A(n801), .B(n128), .O(n798));
  invx g0735(.A(n800), .O(n799));
  orx  g0736(.A(n96), .B(n801), .O(n800));
  orx  g0737(.A(n803), .B(n802), .O(n801));
  andx g0738(.A(n194), .B(n966), .O(n802));
  andx g0739(.A(n804), .B(n182), .O(n803));
  orx  g0740(.A(n806), .B(n805), .O(n804));
  andx g0741(.A(n962), .B(n922), .O(n805));
  andx g0742(.A(n807), .B(n961), .O(n806));
  invx g0743(.A(n922), .O(n807));
  invx g0744(.A(n809), .O(n808));
  orx  g0745(.A(n811), .B(n810), .O(n809));
  andx g0746(.A(n813), .B(n122), .O(n810));
  invx g0747(.A(n812), .O(n811));
  orx  g0748(.A(n122), .B(n813), .O(n812));
  orx  g0749(.A(n815), .B(n814), .O(n813));
  andx g0750(.A(n899), .B(n978), .O(n814));
  andx g0751(.A(n816), .B(n181), .O(n815));
  orx  g0752(.A(n818), .B(n817), .O(n816));
  andx g0753(.A(n974), .B(n920), .O(n817));
  andx g0754(.A(n819), .B(n973), .O(n818));
  invx g0755(.A(n920), .O(n819));
  invx g0756(.A(n821), .O(n820));
  orx  g0757(.A(n823), .B(n822), .O(n821));
  andx g0758(.A(n825), .B(n90), .O(n822));
  invx g0759(.A(n824), .O(n823));
  orx  g0760(.A(n118), .B(n825), .O(n824));
  orx  g0761(.A(n827), .B(n826), .O(n825));
  andx g0762(.A(n194), .B(n990), .O(n826));
  andx g0763(.A(n828), .B(n182), .O(n827));
  orx  g0764(.A(n830), .B(n829), .O(n828));
  andx g0765(.A(n986), .B(n918), .O(n829));
  andx g0766(.A(n831), .B(n985), .O(n830));
  invx g0767(.A(n918), .O(n831));
  invx g0768(.A(n833), .O(n832));
  orx  g0769(.A(n835), .B(n834), .O(n833));
  andx g0770(.A(n837), .B(n112), .O(n834));
  invx g0771(.A(n836), .O(n835));
  orx  g0772(.A(n113), .B(n837), .O(n836));
  orx  g0773(.A(n839), .B(n838), .O(n837));
  andx g0774(.A(n899), .B(n1002), .O(n838));
  andx g0775(.A(n840), .B(n181), .O(n839));
  orx  g0776(.A(n842), .B(n841), .O(n840));
  andx g0777(.A(n998), .B(n916), .O(n841));
  andx g0778(.A(n843), .B(n997), .O(n842));
  invx g0779(.A(n916), .O(n843));
  invx g0780(.A(n845), .O(n844));
  orx  g0781(.A(n847), .B(n846), .O(n845));
  andx g0782(.A(n849), .B(n214), .O(n846));
  invx g0783(.A(n848), .O(n847));
  orx  g0784(.A(n212), .B(n849), .O(n848));
  orx  g0785(.A(n851), .B(n850), .O(n849));
  andx g0786(.A(n194), .B(n1014), .O(n850));
  andx g0787(.A(n852), .B(n182), .O(n851));
  orx  g0788(.A(n854), .B(n853), .O(n852));
  andx g0789(.A(n1010), .B(n914), .O(n853));
  andx g0790(.A(n855), .B(n1009), .O(n854));
  invx g0791(.A(n914), .O(n855));
  invx g0792(.A(n857), .O(n856));
  orx  g0793(.A(n859), .B(n858), .O(n857));
  andx g0794(.A(n861), .B(n208), .O(n858));
  invx g0795(.A(n860), .O(n859));
  orx  g0796(.A(n208), .B(n861), .O(n860));
  orx  g0797(.A(n863), .B(n862), .O(n861));
  andx g0798(.A(n899), .B(n1026), .O(n862));
  andx g0799(.A(n864), .B(n181), .O(n863));
  orx  g0800(.A(n866), .B(n865), .O(n864));
  andx g0801(.A(n1022), .B(n912), .O(n865));
  andx g0802(.A(n867), .B(n1021), .O(n866));
  invx g0803(.A(n912), .O(n867));
  invx g0804(.A(n869), .O(n868));
  orx  g0805(.A(n871), .B(n870), .O(n869));
  andx g0806(.A(n873), .B(n198), .O(n870));
  invx g0807(.A(n872), .O(n871));
  orx  g0808(.A(n197), .B(n873), .O(n872));
  orx  g0809(.A(n875), .B(n874), .O(n873));
  andx g0810(.A(n194), .B(n1038), .O(n874));
  andx g0811(.A(n876), .B(n182), .O(n875));
  orx  g0812(.A(n878), .B(n877), .O(n876));
  andx g0813(.A(n1034), .B(n910), .O(n877));
  andx g0814(.A(n879), .B(n1033), .O(n878));
  invx g0815(.A(n910), .O(n879));
  invx g0816(.A(n881), .O(n880));
  orx  g0817(.A(n883), .B(n882), .O(n881));
  andx g0818(.A(n885), .B(n143), .O(n882));
  invx g0819(.A(n884), .O(n883));
  orx  g0820(.A(n3527), .B(n885), .O(n884));
  orx  g0821(.A(n887), .B(n886), .O(n885));
  andx g0822(.A(n899), .B(n1050), .O(n886));
  andx g0823(.A(n888), .B(n181), .O(n887));
  orx  g0824(.A(n890), .B(n889), .O(n888));
  andx g0825(.A(n1046), .B(n908), .O(n889));
  andx g0826(.A(n891), .B(n1045), .O(n890));
  invx g0827(.A(n908), .O(n891));
  invx g0828(.A(n893), .O(n892));
  andx g0829(.A(n896), .B(n894), .O(n893));
  invx g0830(.A(n895), .O(n894));
  andx g0831(.A(n897), .B(n141), .O(n895));
  orx  g0832(.A(n3528), .B(n897), .O(n896));
  orx  g0833(.A(n900), .B(n898), .O(n897));
  andx g0834(.A(n194), .B(n1062), .O(n898));
  invx g0835(.A(n181), .O(n899));
  andx g0836(.A(n905), .B(n182), .O(n900));
  orx  g0837(.A(n903), .B(n902), .O(n901));
  andx g0838(.A(n3511), .B(n1062), .O(n902));
  andx g0839(.A(n904), .B(n1058), .O(n903));
  andx g0840(.A(n3512), .B(n906), .O(n904));
  andx g0841(.A(n1057), .B(n906), .O(n905));
  orx  g0842(.A(n907), .B(n1047), .O(n906));
  andx g0843(.A(n1045), .B(n908), .O(n907));
  orx  g0844(.A(n909), .B(n1035), .O(n908));
  andx g0845(.A(n1033), .B(n910), .O(n909));
  orx  g0846(.A(n911), .B(n1023), .O(n910));
  andx g0847(.A(n1021), .B(n912), .O(n911));
  orx  g0848(.A(n913), .B(n1011), .O(n912));
  andx g0849(.A(n1009), .B(n914), .O(n913));
  orx  g0850(.A(n915), .B(n999), .O(n914));
  andx g0851(.A(n997), .B(n916), .O(n915));
  orx  g0852(.A(n917), .B(n987), .O(n916));
  andx g0853(.A(n985), .B(n918), .O(n917));
  orx  g0854(.A(n919), .B(n975), .O(n918));
  andx g0855(.A(n973), .B(n920), .O(n919));
  orx  g0856(.A(n921), .B(n963), .O(n920));
  andx g0857(.A(n961), .B(n922), .O(n921));
  orx  g0858(.A(n923), .B(n951), .O(n922));
  andx g0859(.A(n949), .B(n924), .O(n923));
  orx  g0860(.A(n925), .B(n940), .O(n924));
  andx g0861(.A(n938), .B(n926), .O(n925));
  orx  g0862(.A(n928), .B(n927), .O(n926));
  andx g0863(.A(n934), .B(n217), .O(n927));
  andx g0864(.A(n929), .B(n79), .O(n928));
  invx g0865(.A(n930), .O(n929));
  andx g0866(.A(n932), .B(n931), .O(n930));
  orx  g0867(.A(n934), .B(pi03), .O(n931));
  invx g0868(.A(n933), .O(n932));
  andx g0869(.A(pi03), .B(n934), .O(n933));
  orx  g0870(.A(n936), .B(n935), .O(n934));
  andx g0871(.A(n68), .B(n151), .O(n935));
  andx g0872(.A(pi08), .B(n937), .O(n936));
  orx  g0873(.A(n101), .B(n3500), .O(n937));
  invx g0874(.A(n939), .O(n938));
  orx  g0875(.A(n941), .B(n940), .O(n939));
  andx g0876(.A(n943), .B(n3518), .O(n940));
  invx g0877(.A(n942), .O(n941));
  orx  g0878(.A(n943), .B(n139), .O(n942));
  orx  g0879(.A(n948), .B(n944), .O(n943));
  andx g0880(.A(n945), .B(n150), .O(n944));
  andx g0881(.A(n947), .B(n946), .O(n945));
  orx  g0882(.A(n69), .B(n1091), .O(n946));
  orx  g0883(.A(n68), .B(n1092), .O(n947));
  andx g0884(.A(n102), .B(n1096), .O(n948));
  invx g0885(.A(n950), .O(n949));
  orx  g0886(.A(n952), .B(n951), .O(n950));
  andx g0887(.A(n954), .B(n136), .O(n951));
  invx g0888(.A(n953), .O(n952));
  orx  g0889(.A(n954), .B(n135), .O(n953));
  orx  g0890(.A(n956), .B(n955), .O(n954));
  andx g0891(.A(n101), .B(n1105), .O(n955));
  andx g0892(.A(n957), .B(n151), .O(n956));
  orx  g0893(.A(n959), .B(n958), .O(n957));
  andx g0894(.A(n1101), .B(n1088), .O(n958));
  andx g0895(.A(n960), .B(n1100), .O(n959));
  invx g0896(.A(n1088), .O(n960));
  invx g0897(.A(n962), .O(n961));
  orx  g0898(.A(n964), .B(n963), .O(n962));
  andx g0899(.A(n966), .B(n100), .O(n963));
  invx g0900(.A(n965), .O(n964));
  orx  g0901(.A(n966), .B(n100), .O(n965));
  orx  g0902(.A(n968), .B(n967), .O(n966));
  andx g0903(.A(n102), .B(n1116), .O(n967));
  andx g0904(.A(n969), .B(n151), .O(n968));
  orx  g0905(.A(n971), .B(n970), .O(n969));
  andx g0906(.A(n1112), .B(n1086), .O(n970));
  andx g0907(.A(n972), .B(n1111), .O(n971));
  invx g0908(.A(n1086), .O(n972));
  invx g0909(.A(n974), .O(n973));
  orx  g0910(.A(n976), .B(n975), .O(n974));
  andx g0911(.A(n978), .B(n95), .O(n975));
  invx g0912(.A(n977), .O(n976));
  orx  g0913(.A(n73), .B(n978), .O(n977));
  orx  g0914(.A(n980), .B(n979), .O(n978));
  andx g0915(.A(n101), .B(n1128), .O(n979));
  andx g0916(.A(n981), .B(n151), .O(n980));
  orx  g0917(.A(n983), .B(n982), .O(n981));
  andx g0918(.A(n1124), .B(n1084), .O(n982));
  andx g0919(.A(n984), .B(n1123), .O(n983));
  invx g0920(.A(n1084), .O(n984));
  invx g0921(.A(n986), .O(n985));
  orx  g0922(.A(n988), .B(n987), .O(n986));
  andx g0923(.A(n990), .B(n94), .O(n987));
  invx g0924(.A(n989), .O(n988));
  orx  g0925(.A(n121), .B(n990), .O(n989));
  orx  g0926(.A(n992), .B(n991), .O(n990));
  andx g0927(.A(n102), .B(n1140), .O(n991));
  andx g0928(.A(n993), .B(n150), .O(n992));
  orx  g0929(.A(n995), .B(n994), .O(n993));
  andx g0930(.A(n1136), .B(n1082), .O(n994));
  andx g0931(.A(n996), .B(n1135), .O(n995));
  invx g0932(.A(n1082), .O(n996));
  invx g0933(.A(n998), .O(n997));
  orx  g0934(.A(n1000), .B(n999), .O(n998));
  andx g0935(.A(n1002), .B(n117), .O(n999));
  invx g0936(.A(n1001), .O(n1000));
  orx  g0937(.A(n118), .B(n1002), .O(n1001));
  orx  g0938(.A(n1004), .B(n1003), .O(n1002));
  andx g0939(.A(n101), .B(n1152), .O(n1003));
  andx g0940(.A(n1005), .B(n151), .O(n1004));
  orx  g0941(.A(n1007), .B(n1006), .O(n1005));
  andx g0942(.A(n1148), .B(n1080), .O(n1006));
  andx g0943(.A(n1008), .B(n1147), .O(n1007));
  invx g0944(.A(n1080), .O(n1008));
  invx g0945(.A(n1010), .O(n1009));
  orx  g0946(.A(n1012), .B(n1011), .O(n1010));
  andx g0947(.A(n1014), .B(n112), .O(n1011));
  invx g0948(.A(n1013), .O(n1012));
  orx  g0949(.A(n112), .B(n1014), .O(n1013));
  orx  g0950(.A(n1016), .B(n1015), .O(n1014));
  andx g0951(.A(n102), .B(n1164), .O(n1015));
  andx g0952(.A(n1017), .B(n1065), .O(n1016));
  orx  g0953(.A(n1019), .B(n1018), .O(n1017));
  andx g0954(.A(n1160), .B(n1078), .O(n1018));
  andx g0955(.A(n1020), .B(n1159), .O(n1019));
  invx g0956(.A(n1078), .O(n1020));
  invx g0957(.A(n1022), .O(n1021));
  orx  g0958(.A(n1024), .B(n1023), .O(n1022));
  andx g0959(.A(n1026), .B(n213), .O(n1023));
  invx g0960(.A(n1025), .O(n1024));
  orx  g0961(.A(n215), .B(n1026), .O(n1025));
  orx  g0962(.A(n1028), .B(n1027), .O(n1026));
  andx g0963(.A(n101), .B(n1176), .O(n1027));
  andx g0964(.A(n1029), .B(n151), .O(n1028));
  orx  g0965(.A(n1031), .B(n1030), .O(n1029));
  andx g0966(.A(n1172), .B(n1076), .O(n1030));
  andx g0967(.A(n1032), .B(n1171), .O(n1031));
  invx g0968(.A(n1076), .O(n1032));
  invx g0969(.A(n1034), .O(n1033));
  orx  g0970(.A(n1036), .B(n1035), .O(n1034));
  andx g0971(.A(n1038), .B(n211), .O(n1035));
  invx g0972(.A(n1037), .O(n1036));
  orx  g0973(.A(n211), .B(n1038), .O(n1037));
  orx  g0974(.A(n1040), .B(n1039), .O(n1038));
  andx g0975(.A(n102), .B(n1188), .O(n1039));
  andx g0976(.A(n1041), .B(n150), .O(n1040));
  orx  g0977(.A(n1043), .B(n1042), .O(n1041));
  andx g0978(.A(n1184), .B(n1074), .O(n1042));
  andx g0979(.A(n1044), .B(n1183), .O(n1043));
  invx g0980(.A(n1074), .O(n1044));
  invx g0981(.A(n1046), .O(n1045));
  orx  g0982(.A(n1048), .B(n1047), .O(n1046));
  andx g0983(.A(n1050), .B(n197), .O(n1047));
  invx g0984(.A(n1049), .O(n1048));
  orx  g0985(.A(n199), .B(n1050), .O(n1049));
  orx  g0986(.A(n1052), .B(n1051), .O(n1050));
  andx g0987(.A(n101), .B(n1200), .O(n1051));
  andx g0988(.A(n1053), .B(n150), .O(n1052));
  orx  g0989(.A(n1055), .B(n1054), .O(n1053));
  andx g0990(.A(n1196), .B(n1072), .O(n1054));
  andx g0991(.A(n1056), .B(n1195), .O(n1055));
  invx g0992(.A(n1072), .O(n1056));
  invx g0993(.A(n1058), .O(n1057));
  andx g0994(.A(n1061), .B(n1059), .O(n1058));
  invx g0995(.A(n1060), .O(n1059));
  andx g0996(.A(n1062), .B(n144), .O(n1060));
  orx  g0997(.A(n143), .B(n1062), .O(n1061));
  orx  g0998(.A(n1064), .B(n1063), .O(n1062));
  andx g0999(.A(n102), .B(n1212), .O(n1063));
  andx g1000(.A(n1069), .B(n150), .O(n1064));
  orx  g1001(.A(n1067), .B(n1066), .O(n1065));
  andx g1002(.A(n3510), .B(n1212), .O(n1066));
  andx g1003(.A(n1068), .B(n1208), .O(n1067));
  andx g1004(.A(n3511), .B(n1070), .O(n1068));
  andx g1005(.A(n1207), .B(n1070), .O(n1069));
  orx  g1006(.A(n1071), .B(n1197), .O(n1070));
  andx g1007(.A(n1195), .B(n1072), .O(n1071));
  orx  g1008(.A(n1073), .B(n1185), .O(n1072));
  andx g1009(.A(n1183), .B(n1074), .O(n1073));
  orx  g1010(.A(n1075), .B(n1173), .O(n1074));
  andx g1011(.A(n1171), .B(n1076), .O(n1075));
  orx  g1012(.A(n1077), .B(n1161), .O(n1076));
  andx g1013(.A(n1159), .B(n1078), .O(n1077));
  orx  g1014(.A(n1079), .B(n1149), .O(n1078));
  andx g1015(.A(n1147), .B(n1080), .O(n1079));
  orx  g1016(.A(n1081), .B(n1137), .O(n1080));
  andx g1017(.A(n1135), .B(n1082), .O(n1081));
  orx  g1018(.A(n1083), .B(n1125), .O(n1082));
  andx g1019(.A(n1123), .B(n1084), .O(n1083));
  orx  g1020(.A(n1085), .B(n1113), .O(n1084));
  andx g1021(.A(n1111), .B(n1086), .O(n1085));
  orx  g1022(.A(n1087), .B(n1102), .O(n1086));
  andx g1023(.A(n1100), .B(n1088), .O(n1087));
  orx  g1024(.A(n1090), .B(n1089), .O(n1088));
  andx g1025(.A(n1096), .B(n216), .O(n1089));
  andx g1026(.A(n1091), .B(n69), .O(n1090));
  invx g1027(.A(n1092), .O(n1091));
  andx g1028(.A(n1094), .B(n1093), .O(n1092));
  orx  g1029(.A(n1096), .B(pi03), .O(n1093));
  invx g1030(.A(n1095), .O(n1094));
  andx g1031(.A(pi03), .B(n1096), .O(n1095));
  orx  g1032(.A(n1098), .B(n1097), .O(n1096));
  andx g1033(.A(n88), .B(n146), .O(n1097));
  andx g1034(.A(pi10), .B(n1099), .O(n1098));
  orx  g1035(.A(n97), .B(n126), .O(n1099));
  invx g1036(.A(n1101), .O(n1100));
  orx  g1037(.A(n1103), .B(n1102), .O(n1101));
  andx g1038(.A(n1105), .B(n139), .O(n1102));
  invx g1039(.A(n1104), .O(n1103));
  orx  g1040(.A(n1105), .B(n71), .O(n1104));
  orx  g1041(.A(n1110), .B(n1106), .O(n1105));
  andx g1042(.A(n1107), .B(n145), .O(n1106));
  andx g1043(.A(n1109), .B(n1108), .O(n1107));
  orx  g1044(.A(n89), .B(n1239), .O(n1108));
  orx  g1045(.A(n88), .B(n1240), .O(n1109));
  andx g1046(.A(n97), .B(n1244), .O(n1110));
  invx g1047(.A(n1112), .O(n1111));
  orx  g1048(.A(n1114), .B(n1113), .O(n1112));
  andx g1049(.A(n1116), .B(n134), .O(n1113));
  invx g1050(.A(n1115), .O(n1114));
  orx  g1051(.A(n1116), .B(n135), .O(n1115));
  orx  g1052(.A(n1118), .B(n1117), .O(n1116));
  andx g1053(.A(n98), .B(n1253), .O(n1117));
  andx g1054(.A(n1119), .B(n145), .O(n1118));
  orx  g1055(.A(n1121), .B(n1120), .O(n1119));
  andx g1056(.A(n1249), .B(n1236), .O(n1120));
  andx g1057(.A(n1122), .B(n1248), .O(n1121));
  invx g1058(.A(n1236), .O(n1122));
  invx g1059(.A(n1124), .O(n1123));
  orx  g1060(.A(n1126), .B(n1125), .O(n1124));
  andx g1061(.A(n1128), .B(n100), .O(n1125));
  invx g1062(.A(n1127), .O(n1126));
  orx  g1063(.A(n1128), .B(n100), .O(n1127));
  orx  g1064(.A(n1130), .B(n1129), .O(n1128));
  andx g1065(.A(n97), .B(n1264), .O(n1129));
  andx g1066(.A(n1131), .B(n145), .O(n1130));
  orx  g1067(.A(n1133), .B(n1132), .O(n1131));
  andx g1068(.A(n1260), .B(n1234), .O(n1132));
  andx g1069(.A(n1134), .B(n1259), .O(n1133));
  invx g1070(.A(n1234), .O(n1134));
  invx g1071(.A(n1136), .O(n1135));
  orx  g1072(.A(n1138), .B(n1137), .O(n1136));
  andx g1073(.A(n1140), .B(n95), .O(n1137));
  invx g1074(.A(n1139), .O(n1138));
  orx  g1075(.A(n96), .B(n1140), .O(n1139));
  orx  g1076(.A(n1142), .B(n1141), .O(n1140));
  andx g1077(.A(n98), .B(n1276), .O(n1141));
  andx g1078(.A(n1143), .B(n146), .O(n1142));
  orx  g1079(.A(n1145), .B(n1144), .O(n1143));
  andx g1080(.A(n1272), .B(n1232), .O(n1144));
  andx g1081(.A(n1146), .B(n1271), .O(n1145));
  invx g1082(.A(n1232), .O(n1146));
  invx g1083(.A(n1148), .O(n1147));
  orx  g1084(.A(n1150), .B(n1149), .O(n1148));
  andx g1085(.A(n1152), .B(n122), .O(n1149));
  invx g1086(.A(n1151), .O(n1150));
  orx  g1087(.A(n3516), .B(n1152), .O(n1151));
  orx  g1088(.A(n1154), .B(n1153), .O(n1152));
  andx g1089(.A(n97), .B(n1288), .O(n1153));
  andx g1090(.A(n1155), .B(n145), .O(n1154));
  orx  g1091(.A(n1157), .B(n1156), .O(n1155));
  andx g1092(.A(n1284), .B(n1230), .O(n1156));
  andx g1093(.A(n1158), .B(n1283), .O(n1157));
  invx g1094(.A(n1230), .O(n1158));
  invx g1095(.A(n1160), .O(n1159));
  orx  g1096(.A(n1162), .B(n1161), .O(n1160));
  andx g1097(.A(n1164), .B(n118), .O(n1161));
  invx g1098(.A(n1163), .O(n1162));
  orx  g1099(.A(n3523), .B(n1164), .O(n1163));
  orx  g1100(.A(n1166), .B(n1165), .O(n1164));
  andx g1101(.A(n98), .B(n1300), .O(n1165));
  andx g1102(.A(n1167), .B(n146), .O(n1166));
  orx  g1103(.A(n1169), .B(n1168), .O(n1167));
  andx g1104(.A(n1296), .B(n1228), .O(n1168));
  andx g1105(.A(n1170), .B(n1295), .O(n1169));
  invx g1106(.A(n1228), .O(n1170));
  invx g1107(.A(n1172), .O(n1171));
  orx  g1108(.A(n1174), .B(n1173), .O(n1172));
  andx g1109(.A(n1176), .B(n3524), .O(n1173));
  invx g1110(.A(n1175), .O(n1174));
  orx  g1111(.A(n3524), .B(n1176), .O(n1175));
  orx  g1112(.A(n1178), .B(n1177), .O(n1176));
  andx g1113(.A(n97), .B(n1312), .O(n1177));
  andx g1114(.A(n1179), .B(n146), .O(n1178));
  orx  g1115(.A(n1181), .B(n1180), .O(n1179));
  andx g1116(.A(n1308), .B(n1226), .O(n1180));
  andx g1117(.A(n1182), .B(n1307), .O(n1181));
  invx g1118(.A(n1226), .O(n1182));
  invx g1119(.A(n1184), .O(n1183));
  orx  g1120(.A(n1186), .B(n1185), .O(n1184));
  andx g1121(.A(n1188), .B(n212), .O(n1185));
  invx g1122(.A(n1187), .O(n1186));
  orx  g1123(.A(n214), .B(n1188), .O(n1187));
  orx  g1124(.A(n1190), .B(n1189), .O(n1188));
  andx g1125(.A(n98), .B(n1324), .O(n1189));
  andx g1126(.A(n1191), .B(n146), .O(n1190));
  orx  g1127(.A(n1193), .B(n1192), .O(n1191));
  andx g1128(.A(n1320), .B(n1224), .O(n1192));
  andx g1129(.A(n1194), .B(n1319), .O(n1193));
  invx g1130(.A(n1224), .O(n1194));
  invx g1131(.A(n1196), .O(n1195));
  orx  g1132(.A(n1198), .B(n1197), .O(n1196));
  andx g1133(.A(n1200), .B(n210), .O(n1197));
  invx g1134(.A(n1199), .O(n1198));
  orx  g1135(.A(n210), .B(n1200), .O(n1199));
  orx  g1136(.A(n1202), .B(n1201), .O(n1200));
  andx g1137(.A(n97), .B(n1336), .O(n1201));
  andx g1138(.A(n1203), .B(n145), .O(n1202));
  orx  g1139(.A(n1205), .B(n1204), .O(n1203));
  andx g1140(.A(n1332), .B(n1222), .O(n1204));
  andx g1141(.A(n1206), .B(n1331), .O(n1205));
  invx g1142(.A(n1222), .O(n1206));
  invx g1143(.A(n1208), .O(n1207));
  andx g1144(.A(n1211), .B(n1209), .O(n1208));
  invx g1145(.A(n1210), .O(n1209));
  andx g1146(.A(n1212), .B(n199), .O(n1210));
  orx  g1147(.A(n198), .B(n1212), .O(n1211));
  orx  g1148(.A(n1214), .B(n1213), .O(n1212));
  andx g1149(.A(n98), .B(n1348), .O(n1213));
  andx g1150(.A(n1219), .B(n1215), .O(n1214));
  orx  g1151(.A(n1217), .B(n1216), .O(n1215));
  andx g1152(.A(n3509), .B(n1348), .O(n1216));
  andx g1153(.A(n1218), .B(n1344), .O(n1217));
  andx g1154(.A(n3510), .B(n1220), .O(n1218));
  andx g1155(.A(n1343), .B(n1220), .O(n1219));
  orx  g1156(.A(n1221), .B(n1333), .O(n1220));
  andx g1157(.A(n1331), .B(n1222), .O(n1221));
  orx  g1158(.A(n1223), .B(n1321), .O(n1222));
  andx g1159(.A(n1319), .B(n1224), .O(n1223));
  orx  g1160(.A(n1225), .B(n1309), .O(n1224));
  andx g1161(.A(n1307), .B(n1226), .O(n1225));
  orx  g1162(.A(n1227), .B(n1297), .O(n1226));
  andx g1163(.A(n1295), .B(n1228), .O(n1227));
  orx  g1164(.A(n1229), .B(n1285), .O(n1228));
  andx g1165(.A(n1283), .B(n1230), .O(n1229));
  orx  g1166(.A(n1231), .B(n1273), .O(n1230));
  andx g1167(.A(n1271), .B(n1232), .O(n1231));
  orx  g1168(.A(n1233), .B(n1261), .O(n1232));
  andx g1169(.A(n1259), .B(n1234), .O(n1233));
  orx  g1170(.A(n1235), .B(n1250), .O(n1234));
  andx g1171(.A(n1248), .B(n1236), .O(n1235));
  orx  g1172(.A(n1238), .B(n1237), .O(n1236));
  andx g1173(.A(n1244), .B(n164), .O(n1237));
  andx g1174(.A(n1239), .B(n89), .O(n1238));
  invx g1175(.A(n1240), .O(n1239));
  andx g1176(.A(n1242), .B(n1241), .O(n1240));
  orx  g1177(.A(n1244), .B(pi03), .O(n1241));
  invx g1178(.A(n1243), .O(n1242));
  andx g1179(.A(pi03), .B(n1244), .O(n1243));
  orx  g1180(.A(n1246), .B(n1245), .O(n1244));
  andx g1181(.A(n64), .B(n192), .O(n1245));
  andx g1182(.A(pi12), .B(n1247), .O(n1246));
  orx  g1183(.A(n123), .B(n175), .O(n1247));
  invx g1184(.A(n1249), .O(n1248));
  orx  g1185(.A(n1251), .B(n1250), .O(n1249));
  andx g1186(.A(n1253), .B(n108), .O(n1250));
  invx g1187(.A(n1252), .O(n1251));
  orx  g1188(.A(n1253), .B(n108), .O(n1252));
  orx  g1189(.A(n1258), .B(n1254), .O(n1253));
  andx g1190(.A(n1255), .B(n192), .O(n1254));
  andx g1191(.A(n1257), .B(n1256), .O(n1255));
  orx  g1192(.A(n65), .B(n1377), .O(n1256));
  orx  g1193(.A(n64), .B(n1378), .O(n1257));
  andx g1194(.A(n1382), .B(n176), .O(n1258));
  invx g1195(.A(n1260), .O(n1259));
  orx  g1196(.A(n1262), .B(n1261), .O(n1260));
  andx g1197(.A(n1264), .B(n3517), .O(n1261));
  invx g1198(.A(n1263), .O(n1262));
  orx  g1199(.A(n1264), .B(n3517), .O(n1263));
  orx  g1200(.A(n1270), .B(n1265), .O(n1264));
  andx g1201(.A(n1266), .B(n192), .O(n1265));
  orx  g1202(.A(n1268), .B(n1267), .O(n1266));
  andx g1203(.A(n1387), .B(n1374), .O(n1267));
  andx g1204(.A(n1269), .B(n1386), .O(n1268));
  invx g1205(.A(n1374), .O(n1269));
  andx g1206(.A(n1391), .B(n175), .O(n1270));
  invx g1207(.A(n1272), .O(n1271));
  orx  g1208(.A(n1274), .B(n1273), .O(n1272));
  andx g1209(.A(n1276), .B(n100), .O(n1273));
  invx g1210(.A(n1275), .O(n1274));
  orx  g1211(.A(n1276), .B(n100), .O(n1275));
  orx  g1212(.A(n1282), .B(n1277), .O(n1276));
  andx g1213(.A(n1278), .B(n1350), .O(n1277));
  orx  g1214(.A(n1280), .B(n1279), .O(n1278));
  andx g1215(.A(n1398), .B(n1372), .O(n1279));
  andx g1216(.A(n1281), .B(n1397), .O(n1280));
  invx g1217(.A(n1372), .O(n1281));
  andx g1218(.A(n1402), .B(n176), .O(n1282));
  invx g1219(.A(n1284), .O(n1283));
  orx  g1220(.A(n1286), .B(n1285), .O(n1284));
  andx g1221(.A(n1288), .B(n127), .O(n1285));
  invx g1222(.A(n1287), .O(n1286));
  orx  g1223(.A(n127), .B(n1288), .O(n1287));
  orx  g1224(.A(n1294), .B(n1289), .O(n1288));
  andx g1225(.A(n1290), .B(n192), .O(n1289));
  orx  g1226(.A(n1292), .B(n1291), .O(n1290));
  andx g1227(.A(n1410), .B(n1370), .O(n1291));
  andx g1228(.A(n1293), .B(n1409), .O(n1292));
  invx g1229(.A(n1370), .O(n1293));
  andx g1230(.A(n1414), .B(n175), .O(n1294));
  invx g1231(.A(n1296), .O(n1295));
  orx  g1232(.A(n1298), .B(n1297), .O(n1296));
  andx g1233(.A(n1300), .B(n72), .O(n1297));
  invx g1234(.A(n1299), .O(n1298));
  orx  g1235(.A(n72), .B(n1300), .O(n1299));
  orx  g1236(.A(n1306), .B(n1301), .O(n1300));
  andx g1237(.A(n1302), .B(n1350), .O(n1301));
  orx  g1238(.A(n1304), .B(n1303), .O(n1302));
  andx g1239(.A(n1422), .B(n1368), .O(n1303));
  andx g1240(.A(n1305), .B(n1421), .O(n1304));
  invx g1241(.A(n1368), .O(n1305));
  andx g1242(.A(n1426), .B(n176), .O(n1306));
  invx g1243(.A(n1308), .O(n1307));
  orx  g1244(.A(n1310), .B(n1309), .O(n1308));
  andx g1245(.A(n1312), .B(n119), .O(n1309));
  invx g1246(.A(n1311), .O(n1310));
  orx  g1247(.A(n116), .B(n1312), .O(n1311));
  orx  g1248(.A(n1318), .B(n1313), .O(n1312));
  andx g1249(.A(n1314), .B(n192), .O(n1313));
  orx  g1250(.A(n1316), .B(n1315), .O(n1314));
  andx g1251(.A(n1434), .B(n1366), .O(n1315));
  andx g1252(.A(n1317), .B(n1433), .O(n1316));
  invx g1253(.A(n1366), .O(n1317));
  andx g1254(.A(n1438), .B(n175), .O(n1318));
  invx g1255(.A(n1320), .O(n1319));
  orx  g1256(.A(n1322), .B(n1321), .O(n1320));
  andx g1257(.A(n1324), .B(n114), .O(n1321));
  invx g1258(.A(n1323), .O(n1322));
  orx  g1259(.A(n112), .B(n1324), .O(n1323));
  orx  g1260(.A(n1330), .B(n1325), .O(n1324));
  andx g1261(.A(n1326), .B(n1350), .O(n1325));
  orx  g1262(.A(n1328), .B(n1327), .O(n1326));
  andx g1263(.A(n1446), .B(n1364), .O(n1327));
  andx g1264(.A(n1329), .B(n1445), .O(n1328));
  invx g1265(.A(n1364), .O(n1329));
  andx g1266(.A(n1450), .B(n176), .O(n1330));
  invx g1267(.A(n1332), .O(n1331));
  orx  g1268(.A(n1334), .B(n1333), .O(n1332));
  andx g1269(.A(n1336), .B(n215), .O(n1333));
  invx g1270(.A(n1335), .O(n1334));
  orx  g1271(.A(n213), .B(n1336), .O(n1335));
  orx  g1272(.A(n1342), .B(n1337), .O(n1336));
  andx g1273(.A(n1338), .B(n192), .O(n1337));
  orx  g1274(.A(n1340), .B(n1339), .O(n1338));
  andx g1275(.A(n1458), .B(n1362), .O(n1339));
  andx g1276(.A(n1341), .B(n1457), .O(n1340));
  invx g1277(.A(n1362), .O(n1341));
  andx g1278(.A(n1462), .B(n175), .O(n1342));
  invx g1279(.A(n1344), .O(n1343));
  andx g1280(.A(n1347), .B(n1345), .O(n1344));
  invx g1281(.A(n1346), .O(n1345));
  andx g1282(.A(n1348), .B(n209), .O(n1346));
  orx  g1283(.A(n209), .B(n1348), .O(n1347));
  orx  g1284(.A(n1352), .B(n1349), .O(n1348));
  andx g1285(.A(n1351), .B(n1350), .O(n1349));
  invx g1286(.A(n175), .O(n1350));
  andx g1287(.A(n1356), .B(n1360), .O(n1351));
  andx g1288(.A(n1471), .B(n176), .O(n1352));
  orx  g1289(.A(n1354), .B(n2906), .O(n1353));
  andx g1290(.A(n1469), .B(n1355), .O(n1354));
  orx  g1291(.A(n1359), .B(n1356), .O(n1355));
  orx  g1292(.A(n1358), .B(n1357), .O(n1356));
  andx g1293(.A(n1471), .B(n214), .O(n1357));
  andx g1294(.A(pi19), .B(n1470), .O(n1358));
  invx g1295(.A(n1360), .O(n1359));
  orx  g1296(.A(n1361), .B(n1459), .O(n1360));
  andx g1297(.A(n1457), .B(n1362), .O(n1361));
  orx  g1298(.A(n1363), .B(n1447), .O(n1362));
  andx g1299(.A(n1445), .B(n1364), .O(n1363));
  orx  g1300(.A(n1365), .B(n1435), .O(n1364));
  andx g1301(.A(n1433), .B(n1366), .O(n1365));
  orx  g1302(.A(n1367), .B(n1423), .O(n1366));
  andx g1303(.A(n1421), .B(n1368), .O(n1367));
  orx  g1304(.A(n1369), .B(n1411), .O(n1368));
  andx g1305(.A(n1409), .B(n1370), .O(n1369));
  orx  g1306(.A(n1371), .B(n1399), .O(n1370));
  andx g1307(.A(n1397), .B(n1372), .O(n1371));
  orx  g1308(.A(n1373), .B(n1388), .O(n1372));
  andx g1309(.A(n1386), .B(n1374), .O(n1373));
  orx  g1310(.A(n1376), .B(n1375), .O(n1374));
  andx g1311(.A(n1382), .B(n218), .O(n1375));
  andx g1312(.A(n1377), .B(n65), .O(n1376));
  invx g1313(.A(n1378), .O(n1377));
  andx g1314(.A(n1380), .B(n1379), .O(n1378));
  orx  g1315(.A(n1382), .B(pi03), .O(n1379));
  invx g1316(.A(n1381), .O(n1380));
  andx g1317(.A(pi03), .B(n1382), .O(n1381));
  orx  g1318(.A(n1384), .B(n1383), .O(n1382));
  andx g1319(.A(n80), .B(n156), .O(n1383));
  andx g1320(.A(pi14), .B(n1385), .O(n1384));
  orx  g1321(.A(n1473), .B(n126), .O(n1385));
  invx g1322(.A(n1387), .O(n1386));
  orx  g1323(.A(n1389), .B(n1388), .O(n1387));
  andx g1324(.A(n1391), .B(n137), .O(n1388));
  invx g1325(.A(n1390), .O(n1389));
  orx  g1326(.A(n1391), .B(n71), .O(n1390));
  orx  g1327(.A(n1396), .B(n1392), .O(n1391));
  andx g1328(.A(n1393), .B(n155), .O(n1392));
  andx g1329(.A(n1395), .B(n1394), .O(n1393));
  orx  g1330(.A(n81), .B(n1495), .O(n1394));
  orx  g1331(.A(n80), .B(n1496), .O(n1395));
  andx g1332(.A(n188), .B(n1500), .O(n1396));
  invx g1333(.A(n1398), .O(n1397));
  orx  g1334(.A(n1400), .B(n1399), .O(n1398));
  andx g1335(.A(n1402), .B(n134), .O(n1399));
  invx g1336(.A(n1401), .O(n1400));
  orx  g1337(.A(n1402), .B(n134), .O(n1401));
  orx  g1338(.A(n1404), .B(n1403), .O(n1402));
  andx g1339(.A(n188), .B(n1509), .O(n1403));
  andx g1340(.A(n1405), .B(n156), .O(n1404));
  orx  g1341(.A(n1407), .B(n1406), .O(n1405));
  andx g1342(.A(n1505), .B(n1492), .O(n1406));
  andx g1343(.A(n1408), .B(n1504), .O(n1407));
  invx g1344(.A(n1492), .O(n1408));
  invx g1345(.A(n1410), .O(n1409));
  orx  g1346(.A(n1412), .B(n1411), .O(n1410));
  andx g1347(.A(n1414), .B(n100), .O(n1411));
  invx g1348(.A(n1413), .O(n1412));
  orx  g1349(.A(n1414), .B(n100), .O(n1413));
  orx  g1350(.A(n1416), .B(n1415), .O(n1414));
  andx g1351(.A(n188), .B(n1520), .O(n1415));
  andx g1352(.A(n1417), .B(n155), .O(n1416));
  orx  g1353(.A(n1419), .B(n1418), .O(n1417));
  andx g1354(.A(n1516), .B(n1490), .O(n1418));
  andx g1355(.A(n1420), .B(n1515), .O(n1419));
  invx g1356(.A(n1490), .O(n1420));
  invx g1357(.A(n1422), .O(n1421));
  orx  g1358(.A(n1424), .B(n1423), .O(n1422));
  andx g1359(.A(n1426), .B(n96), .O(n1423));
  invx g1360(.A(n1425), .O(n1424));
  orx  g1361(.A(n128), .B(n1426), .O(n1425));
  orx  g1362(.A(n1428), .B(n1427), .O(n1426));
  andx g1363(.A(n188), .B(n1532), .O(n1427));
  andx g1364(.A(n1429), .B(n156), .O(n1428));
  orx  g1365(.A(n1431), .B(n1430), .O(n1429));
  andx g1366(.A(n1528), .B(n1488), .O(n1430));
  andx g1367(.A(n1432), .B(n1527), .O(n1431));
  invx g1368(.A(n1488), .O(n1432));
  invx g1369(.A(n1434), .O(n1433));
  orx  g1370(.A(n1436), .B(n1435), .O(n1434));
  andx g1371(.A(n1438), .B(n3516), .O(n1435));
  invx g1372(.A(n1437), .O(n1436));
  orx  g1373(.A(n121), .B(n1438), .O(n1437));
  orx  g1374(.A(n1440), .B(n1439), .O(n1438));
  andx g1375(.A(n188), .B(n1544), .O(n1439));
  andx g1376(.A(n1441), .B(n155), .O(n1440));
  orx  g1377(.A(n1443), .B(n1442), .O(n1441));
  andx g1378(.A(n1540), .B(n1486), .O(n1442));
  andx g1379(.A(n1444), .B(n1539), .O(n1443));
  invx g1380(.A(n1486), .O(n1444));
  invx g1381(.A(n1446), .O(n1445));
  orx  g1382(.A(n1448), .B(n1447), .O(n1446));
  andx g1383(.A(n1450), .B(n3523), .O(n1447));
  invx g1384(.A(n1449), .O(n1448));
  orx  g1385(.A(n116), .B(n1450), .O(n1449));
  orx  g1386(.A(n1452), .B(n1451), .O(n1450));
  andx g1387(.A(n188), .B(n1556), .O(n1451));
  andx g1388(.A(n1453), .B(n156), .O(n1452));
  orx  g1389(.A(n1455), .B(n1454), .O(n1453));
  andx g1390(.A(n1552), .B(n1484), .O(n1454));
  andx g1391(.A(n1456), .B(n1551), .O(n1455));
  invx g1392(.A(n1484), .O(n1456));
  invx g1393(.A(n1458), .O(n1457));
  orx  g1394(.A(n1460), .B(n1459), .O(n1458));
  andx g1395(.A(n1462), .B(n114), .O(n1459));
  invx g1396(.A(n1461), .O(n1460));
  orx  g1397(.A(n112), .B(n1462), .O(n1461));
  orx  g1398(.A(n1464), .B(n1463), .O(n1462));
  andx g1399(.A(n1473), .B(n1568), .O(n1463));
  andx g1400(.A(n1465), .B(n155), .O(n1464));
  orx  g1401(.A(n1467), .B(n1466), .O(n1465));
  andx g1402(.A(n1564), .B(n1482), .O(n1466));
  andx g1403(.A(n1468), .B(n1563), .O(n1467));
  invx g1404(.A(n1482), .O(n1468));
  orx  g1405(.A(pi19), .B(n1470), .O(n1469));
  invx g1406(.A(n1471), .O(n1470));
  orx  g1407(.A(n1474), .B(n1472), .O(n1471));
  andx g1408(.A(n1473), .B(n1580), .O(n1472));
  invx g1409(.A(n155), .O(n1473));
  andx g1410(.A(n1479), .B(n156), .O(n1474));
  orx  g1411(.A(n1477), .B(n1476), .O(n1475));
  andx g1412(.A(n3507), .B(n1580), .O(n1476));
  andx g1413(.A(n1478), .B(n1576), .O(n1477));
  andx g1414(.A(n3508), .B(n1480), .O(n1478));
  andx g1415(.A(n1575), .B(n1480), .O(n1479));
  orx  g1416(.A(n1481), .B(n1565), .O(n1480));
  andx g1417(.A(n1563), .B(n1482), .O(n1481));
  orx  g1418(.A(n1483), .B(n1553), .O(n1482));
  andx g1419(.A(n1551), .B(n1484), .O(n1483));
  orx  g1420(.A(n1485), .B(n1541), .O(n1484));
  andx g1421(.A(n1539), .B(n1486), .O(n1485));
  orx  g1422(.A(n1487), .B(n1529), .O(n1486));
  andx g1423(.A(n1527), .B(n1488), .O(n1487));
  orx  g1424(.A(n1489), .B(n1517), .O(n1488));
  andx g1425(.A(n1515), .B(n1490), .O(n1489));
  orx  g1426(.A(n1491), .B(n1506), .O(n1490));
  andx g1427(.A(n1504), .B(n1492), .O(n1491));
  orx  g1428(.A(n1494), .B(n1493), .O(n1492));
  andx g1429(.A(n1500), .B(n217), .O(n1493));
  andx g1430(.A(n1495), .B(n81), .O(n1494));
  invx g1431(.A(n1496), .O(n1495));
  andx g1432(.A(n1498), .B(n1497), .O(n1496));
  orx  g1433(.A(n1500), .B(pi03), .O(n1497));
  invx g1434(.A(n1499), .O(n1498));
  andx g1435(.A(pi03), .B(n1500), .O(n1499));
  orx  g1436(.A(n1502), .B(n1501), .O(n1500));
  andx g1437(.A(n82), .B(n142), .O(n1501));
  andx g1438(.A(pi16), .B(n1503), .O(n1502));
  orx  g1439(.A(n1582), .B(n91), .O(n1503));
  invx g1440(.A(n1505), .O(n1504));
  orx  g1441(.A(n1507), .B(n1506), .O(n1505));
  andx g1442(.A(n1509), .B(n71), .O(n1506));
  invx g1443(.A(n1508), .O(n1507));
  orx  g1444(.A(n1509), .B(n71), .O(n1508));
  orx  g1445(.A(n1514), .B(n1510), .O(n1509));
  andx g1446(.A(n1511), .B(n142), .O(n1510));
  andx g1447(.A(n1513), .B(n1512), .O(n1511));
  orx  g1448(.A(n83), .B(n1602), .O(n1512));
  orx  g1449(.A(n82), .B(n1603), .O(n1513));
  andx g1450(.A(n186), .B(n1607), .O(n1514));
  invx g1451(.A(n1516), .O(n1515));
  orx  g1452(.A(n1518), .B(n1517), .O(n1516));
  andx g1453(.A(n1520), .B(n134), .O(n1517));
  invx g1454(.A(n1519), .O(n1518));
  orx  g1455(.A(n1520), .B(n136), .O(n1519));
  orx  g1456(.A(n1522), .B(n1521), .O(n1520));
  andx g1457(.A(n186), .B(n1616), .O(n1521));
  andx g1458(.A(n1523), .B(n142), .O(n1522));
  orx  g1459(.A(n1525), .B(n1524), .O(n1523));
  andx g1460(.A(n1612), .B(n1599), .O(n1524));
  andx g1461(.A(n1526), .B(n1611), .O(n1525));
  invx g1462(.A(n1599), .O(n1526));
  invx g1463(.A(n1528), .O(n1527));
  orx  g1464(.A(n1530), .B(n1529), .O(n1528));
  andx g1465(.A(n1532), .B(n99), .O(n1529));
  invx g1466(.A(n1531), .O(n1530));
  orx  g1467(.A(n1532), .B(n132), .O(n1531));
  orx  g1468(.A(n1534), .B(n1533), .O(n1532));
  andx g1469(.A(n186), .B(n1627), .O(n1533));
  andx g1470(.A(n1535), .B(n142), .O(n1534));
  orx  g1471(.A(n1537), .B(n1536), .O(n1535));
  andx g1472(.A(n1623), .B(n1597), .O(n1536));
  andx g1473(.A(n1538), .B(n1622), .O(n1537));
  invx g1474(.A(n1597), .O(n1538));
  invx g1475(.A(n1540), .O(n1539));
  orx  g1476(.A(n1542), .B(n1541), .O(n1540));
  andx g1477(.A(n1544), .B(n127), .O(n1541));
  invx g1478(.A(n1543), .O(n1542));
  orx  g1479(.A(n128), .B(n1544), .O(n1543));
  orx  g1480(.A(n1546), .B(n1545), .O(n1544));
  andx g1481(.A(n186), .B(n1639), .O(n1545));
  andx g1482(.A(n1547), .B(n142), .O(n1546));
  orx  g1483(.A(n1549), .B(n1548), .O(n1547));
  andx g1484(.A(n1635), .B(n1595), .O(n1548));
  andx g1485(.A(n1550), .B(n1634), .O(n1549));
  invx g1486(.A(n1595), .O(n1550));
  invx g1487(.A(n1552), .O(n1551));
  orx  g1488(.A(n1554), .B(n1553), .O(n1552));
  andx g1489(.A(n1556), .B(n3516), .O(n1553));
  invx g1490(.A(n1555), .O(n1554));
  orx  g1491(.A(n94), .B(n1556), .O(n1555));
  orx  g1492(.A(n1558), .B(n1557), .O(n1556));
  andx g1493(.A(n1582), .B(n1651), .O(n1557));
  andx g1494(.A(n1559), .B(n142), .O(n1558));
  orx  g1495(.A(n1561), .B(n1560), .O(n1559));
  andx g1496(.A(n1647), .B(n1593), .O(n1560));
  andx g1497(.A(n1562), .B(n1646), .O(n1561));
  invx g1498(.A(n1593), .O(n1562));
  invx g1499(.A(n1564), .O(n1563));
  orx  g1500(.A(n1566), .B(n1565), .O(n1564));
  andx g1501(.A(n1568), .B(n119), .O(n1565));
  invx g1502(.A(n1567), .O(n1566));
  orx  g1503(.A(n116), .B(n1568), .O(n1567));
  orx  g1504(.A(n1570), .B(n1569), .O(n1568));
  andx g1505(.A(n1582), .B(n1663), .O(n1569));
  andx g1506(.A(n1571), .B(n1584), .O(n1570));
  orx  g1507(.A(n1573), .B(n1572), .O(n1571));
  andx g1508(.A(n1659), .B(n1591), .O(n1572));
  andx g1509(.A(n1574), .B(n1658), .O(n1573));
  invx g1510(.A(n1591), .O(n1574));
  invx g1511(.A(n1576), .O(n1575));
  andx g1512(.A(n1579), .B(n1577), .O(n1576));
  invx g1513(.A(n1578), .O(n1577));
  andx g1514(.A(n1580), .B(n114), .O(n1578));
  orx  g1515(.A(n114), .B(n1580), .O(n1579));
  orx  g1516(.A(n1583), .B(n1581), .O(n1580));
  andx g1517(.A(n1582), .B(n1675), .O(n1581));
  invx g1518(.A(n1584), .O(n1582));
  andx g1519(.A(n1588), .B(n1584), .O(n1583));
  orx  g1520(.A(n1586), .B(n1585), .O(n1584));
  andx g1521(.A(n3506), .B(n1675), .O(n1585));
  andx g1522(.A(n1587), .B(n1671), .O(n1586));
  andx g1523(.A(n3507), .B(n1589), .O(n1587));
  andx g1524(.A(n1670), .B(n1589), .O(n1588));
  orx  g1525(.A(n1590), .B(n1660), .O(n1589));
  andx g1526(.A(n1658), .B(n1591), .O(n1590));
  orx  g1527(.A(n1592), .B(n1648), .O(n1591));
  andx g1528(.A(n1646), .B(n1593), .O(n1592));
  orx  g1529(.A(n1594), .B(n1636), .O(n1593));
  andx g1530(.A(n1634), .B(n1595), .O(n1594));
  orx  g1531(.A(n1596), .B(n1624), .O(n1595));
  andx g1532(.A(n1622), .B(n1597), .O(n1596));
  orx  g1533(.A(n1598), .B(n1613), .O(n1597));
  andx g1534(.A(n1611), .B(n1599), .O(n1598));
  orx  g1535(.A(n1601), .B(n1600), .O(n1599));
  andx g1536(.A(n1607), .B(n216), .O(n1600));
  andx g1537(.A(n1602), .B(n83), .O(n1601));
  invx g1538(.A(n1603), .O(n1602));
  andx g1539(.A(n1605), .B(n1604), .O(n1603));
  orx  g1540(.A(n1607), .B(pi03), .O(n1604));
  invx g1541(.A(n1606), .O(n1605));
  andx g1542(.A(pi03), .B(n1607), .O(n1606));
  orx  g1543(.A(n1609), .B(n1608), .O(n1607));
  andx g1544(.A(n84), .B(n1677), .O(n1608));
  andx g1545(.A(pi18), .B(n1610), .O(n1609));
  orx  g1546(.A(n124), .B(n191), .O(n1610));
  invx g1547(.A(n1612), .O(n1611));
  orx  g1548(.A(n1614), .B(n1613), .O(n1612));
  andx g1549(.A(n1616), .B(n139), .O(n1613));
  invx g1550(.A(n1615), .O(n1614));
  orx  g1551(.A(n1616), .B(n137), .O(n1615));
  orx  g1552(.A(n1621), .B(n1617), .O(n1616));
  andx g1553(.A(n1618), .B(n1677), .O(n1617));
  andx g1554(.A(n1620), .B(n1619), .O(n1618));
  orx  g1555(.A(n85), .B(n1698), .O(n1619));
  orx  g1556(.A(n84), .B(n1699), .O(n1620));
  andx g1557(.A(n1703), .B(n191), .O(n1621));
  invx g1558(.A(n1623), .O(n1622));
  orx  g1559(.A(n1625), .B(n1624), .O(n1623));
  andx g1560(.A(n1627), .B(n134), .O(n1624));
  invx g1561(.A(n1626), .O(n1625));
  orx  g1562(.A(n1627), .B(n136), .O(n1626));
  orx  g1563(.A(n1633), .B(n1628), .O(n1627));
  andx g1564(.A(n1629), .B(n1677), .O(n1628));
  orx  g1565(.A(n1631), .B(n1630), .O(n1629));
  andx g1566(.A(n1708), .B(n1695), .O(n1630));
  andx g1567(.A(n1632), .B(n1707), .O(n1631));
  invx g1568(.A(n1695), .O(n1632));
  andx g1569(.A(n1712), .B(n191), .O(n1633));
  invx g1570(.A(n1635), .O(n1634));
  orx  g1571(.A(n1637), .B(n1636), .O(n1635));
  andx g1572(.A(n1639), .B(n99), .O(n1636));
  invx g1573(.A(n1638), .O(n1637));
  orx  g1574(.A(n1639), .B(n99), .O(n1638));
  orx  g1575(.A(n1645), .B(n1640), .O(n1639));
  andx g1576(.A(n1641), .B(n1677), .O(n1640));
  orx  g1577(.A(n1643), .B(n1642), .O(n1641));
  andx g1578(.A(n1719), .B(n1693), .O(n1642));
  andx g1579(.A(n1644), .B(n1718), .O(n1643));
  invx g1580(.A(n1693), .O(n1644));
  andx g1581(.A(n1723), .B(n191), .O(n1645));
  invx g1582(.A(n1647), .O(n1646));
  orx  g1583(.A(n1649), .B(n1648), .O(n1647));
  andx g1584(.A(n1651), .B(n96), .O(n1648));
  invx g1585(.A(n1650), .O(n1649));
  orx  g1586(.A(n95), .B(n1651), .O(n1650));
  orx  g1587(.A(n1657), .B(n1652), .O(n1651));
  andx g1588(.A(n1653), .B(n1677), .O(n1652));
  orx  g1589(.A(n1655), .B(n1654), .O(n1653));
  andx g1590(.A(n1731), .B(n1691), .O(n1654));
  andx g1591(.A(n1656), .B(n1730), .O(n1655));
  invx g1592(.A(n1691), .O(n1656));
  andx g1593(.A(n1735), .B(n191), .O(n1657));
  invx g1594(.A(n1659), .O(n1658));
  orx  g1595(.A(n1661), .B(n1660), .O(n1659));
  andx g1596(.A(n1663), .B(n120), .O(n1660));
  invx g1597(.A(n1662), .O(n1661));
  orx  g1598(.A(n120), .B(n1663), .O(n1662));
  orx  g1599(.A(n1669), .B(n1664), .O(n1663));
  andx g1600(.A(n1665), .B(n1677), .O(n1664));
  orx  g1601(.A(n1667), .B(n1666), .O(n1665));
  andx g1602(.A(n1742), .B(n1689), .O(n1666));
  andx g1603(.A(n1668), .B(n1741), .O(n1667));
  invx g1604(.A(n1689), .O(n1668));
  andx g1605(.A(n1746), .B(n1680), .O(n1669));
  invx g1606(.A(n1671), .O(n1670));
  andx g1607(.A(n1674), .B(n1672), .O(n1671));
  invx g1608(.A(n1673), .O(n1672));
  andx g1609(.A(n1675), .B(n116), .O(n1673));
  orx  g1610(.A(n90), .B(n1675), .O(n1674));
  orx  g1611(.A(n1679), .B(n1676), .O(n1675));
  andx g1612(.A(n1678), .B(n1677), .O(n1676));
  invx g1613(.A(n1680), .O(n1677));
  andx g1614(.A(n1683), .B(n1687), .O(n1678));
  andx g1615(.A(n1755), .B(n1680), .O(n1679));
  orx  g1616(.A(n1681), .B(n3237), .O(n1680));
  andx g1617(.A(n1753), .B(n1682), .O(n1681));
  orx  g1618(.A(n1686), .B(n1683), .O(n1682));
  orx  g1619(.A(n1685), .B(n1684), .O(n1683));
  andx g1620(.A(n1755), .B(n94), .O(n1684));
  andx g1621(.A(pi13), .B(n1754), .O(n1685));
  invx g1622(.A(n1687), .O(n1686));
  orx  g1623(.A(n1688), .B(n1743), .O(n1687));
  andx g1624(.A(n1741), .B(n1689), .O(n1688));
  orx  g1625(.A(n1690), .B(n1732), .O(n1689));
  andx g1626(.A(n1730), .B(n1691), .O(n1690));
  orx  g1627(.A(n1692), .B(n1720), .O(n1691));
  andx g1628(.A(n1718), .B(n1693), .O(n1692));
  orx  g1629(.A(n1694), .B(n1709), .O(n1693));
  andx g1630(.A(n1707), .B(n1695), .O(n1694));
  orx  g1631(.A(n1697), .B(n1696), .O(n1695));
  andx g1632(.A(n1703), .B(n219), .O(n1696));
  andx g1633(.A(n1698), .B(n85), .O(n1697));
  invx g1634(.A(n1699), .O(n1698));
  andx g1635(.A(n1701), .B(n1700), .O(n1699));
  orx  g1636(.A(n1703), .B(pi03), .O(n1700));
  invx g1637(.A(n1702), .O(n1701));
  andx g1638(.A(pi03), .B(n1703), .O(n1702));
  orx  g1639(.A(n1705), .B(n1704), .O(n1703));
  andx g1640(.A(n86), .B(n165), .O(n1704));
  andx g1641(.A(pi20), .B(n1706), .O(n1705));
  orx  g1642(.A(n1757), .B(n125), .O(n1706));
  invx g1643(.A(n1708), .O(n1707));
  orx  g1644(.A(n1710), .B(n1709), .O(n1708));
  andx g1645(.A(n1712), .B(n107), .O(n1709));
  invx g1646(.A(n1711), .O(n1710));
  orx  g1647(.A(n1712), .B(n107), .O(n1711));
  orx  g1648(.A(n1717), .B(n1713), .O(n1712));
  andx g1649(.A(n1714), .B(n165), .O(n1713));
  andx g1650(.A(n1716), .B(n1715), .O(n1714));
  orx  g1651(.A(n87), .B(n1790), .O(n1715));
  orx  g1652(.A(n86), .B(n1791), .O(n1716));
  andx g1653(.A(n1757), .B(n1795), .O(n1717));
  invx g1654(.A(n1719), .O(n1718));
  orx  g1655(.A(n1721), .B(n1720), .O(n1719));
  andx g1656(.A(n1723), .B(n104), .O(n1720));
  invx g1657(.A(n1722), .O(n1721));
  orx  g1658(.A(n1723), .B(n104), .O(n1722));
  orx  g1659(.A(n1725), .B(n1724), .O(n1723));
  andx g1660(.A(n1757), .B(n1804), .O(n1724));
  andx g1661(.A(n1726), .B(n165), .O(n1725));
  orx  g1662(.A(n1728), .B(n1727), .O(n1726));
  andx g1663(.A(n1800), .B(n1787), .O(n1727));
  andx g1664(.A(n1729), .B(n1799), .O(n1728));
  invx g1665(.A(n1787), .O(n1729));
  invx g1666(.A(n1731), .O(n1730));
  orx  g1667(.A(n1733), .B(n1732), .O(n1731));
  andx g1668(.A(n1735), .B(n99), .O(n1732));
  invx g1669(.A(n1734), .O(n1733));
  orx  g1670(.A(n1735), .B(n99), .O(n1734));
  orx  g1671(.A(n1740), .B(n1736), .O(n1735));
  andx g1672(.A(n1737), .B(n165), .O(n1736));
  andx g1673(.A(n1739), .B(n1738), .O(n1737));
  orx  g1674(.A(n1770), .B(n1785), .O(n1738));
  invx g1675(.A(n1769), .O(n1739));
  andx g1676(.A(n1757), .B(n1774), .O(n1740));
  invx g1677(.A(n1742), .O(n1741));
  orx  g1678(.A(n1744), .B(n1743), .O(n1742));
  andx g1679(.A(n1746), .B(n129), .O(n1743));
  invx g1680(.A(n1745), .O(n1744));
  orx  g1681(.A(n128), .B(n1746), .O(n1745));
  orx  g1682(.A(n1748), .B(n1747), .O(n1746));
  andx g1683(.A(n1757), .B(n1815), .O(n1747));
  andx g1684(.A(n1749), .B(n165), .O(n1748));
  orx  g1685(.A(n1751), .B(n1750), .O(n1749));
  andx g1686(.A(n1811), .B(n1767), .O(n1750));
  andx g1687(.A(n1752), .B(n1810), .O(n1751));
  invx g1688(.A(n1767), .O(n1752));
  orx  g1689(.A(pi13), .B(n1754), .O(n1753));
  invx g1690(.A(n1755), .O(n1754));
  orx  g1691(.A(n1758), .B(n1756), .O(n1755));
  andx g1692(.A(n1757), .B(n1828), .O(n1756));
  invx g1693(.A(n165), .O(n1757));
  andx g1694(.A(n1764), .B(n165), .O(n1758));
  orx  g1695(.A(n1761), .B(n1760), .O(n1759));
  andx g1696(.A(n3504), .B(n1828), .O(n1760));
  andx g1697(.A(n1763), .B(n1762), .O(n1761));
  invx g1698(.A(n1824), .O(n1762));
  andx g1699(.A(n3505), .B(n1765), .O(n1763));
  andx g1700(.A(n1824), .B(n1765), .O(n1764));
  orx  g1701(.A(n1766), .B(n1812), .O(n1765));
  andx g1702(.A(n1810), .B(n1767), .O(n1766));
  orx  g1703(.A(n1769), .B(n1768), .O(n1767));
  andx g1704(.A(n1774), .B(n3517), .O(n1768));
  andx g1705(.A(n1785), .B(n1770), .O(n1769));
  orx  g1706(.A(n1773), .B(n1771), .O(n1770));
  invx g1707(.A(n1772), .O(n1771));
  orx  g1708(.A(n1774), .B(pi07), .O(n1772));
  andx g1709(.A(pi07), .B(n1774), .O(n1773));
  orx  g1710(.A(n1778), .B(n1775), .O(n1774));
  andx g1711(.A(n1859), .B(n1776), .O(n1775));
  orx  g1712(.A(n1830), .B(n1777), .O(n1776));
  andx g1713(.A(n1781), .B(n105), .O(n1777));
  andx g1714(.A(n1779), .B(n1831), .O(n1778));
  andx g1715(.A(n1781), .B(n1780), .O(n1779));
  invx g1716(.A(n1850), .O(n1780));
  orx  g1717(.A(n1782), .B(n1851), .O(n1781));
  andx g1718(.A(n1783), .B(n1857), .O(n1782));
  orx  g1719(.A(pi05), .B(n1784), .O(n1783));
  invx g1720(.A(n1859), .O(n1784));
  orx  g1721(.A(n1786), .B(n1801), .O(n1785));
  andx g1722(.A(n1799), .B(n1787), .O(n1786));
  orx  g1723(.A(n1789), .B(n1788), .O(n1787));
  andx g1724(.A(n1795), .B(n218), .O(n1788));
  andx g1725(.A(n1790), .B(n87), .O(n1789));
  invx g1726(.A(n1791), .O(n1790));
  andx g1727(.A(n1793), .B(n1792), .O(n1791));
  orx  g1728(.A(n1795), .B(pi03), .O(n1792));
  invx g1729(.A(n1794), .O(n1793));
  andx g1730(.A(pi03), .B(n1795), .O(n1794));
  orx  g1731(.A(n1797), .B(n1796), .O(n1795));
  andx g1732(.A(n1831), .B(n3419), .O(n1796));
  andx g1733(.A(pi22), .B(n1798), .O(n1797));
  orx  g1734(.A(n126), .B(n1830), .O(n1798));
  invx g1735(.A(n1800), .O(n1799));
  orx  g1736(.A(n1802), .B(n1801), .O(n1800));
  andx g1737(.A(n1804), .B(n139), .O(n1801));
  invx g1738(.A(n1803), .O(n1802));
  orx  g1739(.A(n1804), .B(n105), .O(n1803));
  orx  g1740(.A(n1808), .B(n1805), .O(n1804));
  andx g1741(.A(n1807), .B(n1806), .O(n1805));
  invx g1742(.A(n1853), .O(n1806));
  andx g1743(.A(n1831), .B(n3367), .O(n1807));
  andx g1744(.A(n1809), .B(n1853), .O(n1808));
  orx  g1745(.A(n1830), .B(n3372), .O(n1809));
  invx g1746(.A(n1811), .O(n1810));
  orx  g1747(.A(n1813), .B(n1812), .O(n1811));
  andx g1748(.A(n1815), .B(n3522), .O(n1812));
  invx g1749(.A(n1814), .O(n1813));
  orx  g1750(.A(n1815), .B(n99), .O(n1814));
  orx  g1751(.A(n1823), .B(n1816), .O(n1815));
  andx g1752(.A(n1817), .B(n1831), .O(n1816));
  andx g1753(.A(n1820), .B(n1818), .O(n1817));
  invx g1754(.A(n1819), .O(n1818));
  andx g1755(.A(n1849), .B(n1821), .O(n1819));
  orx  g1756(.A(n1821), .B(n1849), .O(n1820));
  andx g1757(.A(n1839), .B(n1822), .O(n1821));
  invx g1758(.A(n1837), .O(n1822));
  andx g1759(.A(n1840), .B(n1830), .O(n1823));
  andx g1760(.A(n1826), .B(n1825), .O(n1824));
  orx  g1761(.A(n1828), .B(pi11), .O(n1825));
  invx g1762(.A(n1827), .O(n1826));
  andx g1763(.A(pi11), .B(n1828), .O(n1827));
  orx  g1764(.A(n1835), .B(n1829), .O(n1828));
  andx g1765(.A(n1866), .B(n1830), .O(n1829));
  invx g1766(.A(n1831), .O(n1830));
  andx g1767(.A(n1832), .B(n3504), .O(n1831));
  orx  g1768(.A(n1865), .B(n1833), .O(n1832));
  andx g1769(.A(n1836), .B(n1834), .O(n1833));
  orx  g1770(.A(n99), .B(n1866), .O(n1834));
  andx g1771(.A(n1865), .B(n1836), .O(n1835));
  orx  g1772(.A(n1838), .B(n1837), .O(n1836));
  andx g1773(.A(n3517), .B(n1840), .O(n1837));
  andx g1774(.A(n1849), .B(n1839), .O(n1838));
  orx  g1775(.A(n136), .B(n1840), .O(n1839));
  orx  g1776(.A(n1844), .B(n1841), .O(n1840));
  andx g1777(.A(n1885), .B(n1842), .O(n1841));
  orx  g1778(.A(n1868), .B(n1843), .O(n1842));
  andx g1779(.A(n1845), .B(n138), .O(n1843));
  andx g1780(.A(n1847), .B(n1845), .O(n1844));
  orx  g1781(.A(n1846), .B(n1878), .O(n1845));
  andx g1782(.A(pi05), .B(n1877), .O(n1846));
  invx g1783(.A(n1848), .O(n1847));
  orx  g1784(.A(n1868), .B(n1876), .O(n1848));
  orx  g1785(.A(n1850), .B(n1858), .O(n1849));
  andx g1786(.A(n1857), .B(n1851), .O(n1850));
  orx  g1787(.A(n1852), .B(n3415), .O(n1851));
  andx g1788(.A(n3417), .B(n1853), .O(n1852));
  orx  g1789(.A(n1855), .B(n1854), .O(n1853));
  andx g1790(.A(n3455), .B(n1869), .O(n1854));
  andx g1791(.A(pi24), .B(n1856), .O(n1855));
  orx  g1792(.A(n1868), .B(n125), .O(n1856));
  orx  g1793(.A(n138), .B(n1859), .O(n1857));
  andx g1794(.A(n1859), .B(n108), .O(n1858));
  orx  g1795(.A(n1863), .B(n1860), .O(n1859));
  andx g1796(.A(n1862), .B(n1861), .O(n1860));
  invx g1797(.A(n1880), .O(n1861));
  andx g1798(.A(n3431), .B(n1869), .O(n1862));
  andx g1799(.A(n1864), .B(n1880), .O(n1863));
  orx  g1800(.A(n1868), .B(n3436), .O(n1864));
  andx g1801(.A(n130), .B(n1866), .O(n1865));
  orx  g1802(.A(n1874), .B(n1867), .O(n1866));
  andx g1803(.A(n1868), .B(n1891), .O(n1867));
  invx g1804(.A(n1869), .O(n1868));
  orx  g1805(.A(n1871), .B(n1870), .O(n1869));
  andx g1806(.A(n3502), .B(n1891), .O(n1870));
  andx g1807(.A(n1872), .B(n3503), .O(n1871));
  andx g1808(.A(n1875), .B(n1873), .O(n1872));
  orx  g1809(.A(n1891), .B(n133), .O(n1873));
  andx g1810(.A(n1890), .B(n1875), .O(n1874));
  orx  g1811(.A(n1876), .B(n1884), .O(n1875));
  andx g1812(.A(n1878), .B(n1877), .O(n1876));
  orx  g1813(.A(n138), .B(n1885), .O(n1877));
  orx  g1814(.A(n1879), .B(n3451), .O(n1878));
  andx g1815(.A(n3453), .B(n1880), .O(n1879));
  orx  g1816(.A(n1882), .B(n1881), .O(n1880));
  andx g1817(.A(n3459), .B(n1895), .O(n1881));
  andx g1818(.A(pi26), .B(n1883), .O(n1882));
  orx  g1819(.A(n1894), .B(n3500), .O(n1883));
  andx g1820(.A(n1885), .B(n71), .O(n1884));
  orx  g1821(.A(n1888), .B(n1886), .O(n1885));
  andx g1822(.A(n1887), .B(n1903), .O(n1886));
  andx g1823(.A(n3466), .B(n1895), .O(n1887));
  andx g1824(.A(n1889), .B(n1902), .O(n1888));
  orx  g1825(.A(n3480), .B(n1894), .O(n1889));
  andx g1826(.A(n1891), .B(n103), .O(n1890));
  andx g1827(.A(n1892), .B(n1905), .O(n1891));
  orx  g1828(.A(n1894), .B(n1893), .O(n1892));
  andx g1829(.A(n108), .B(n1900), .O(n1893));
  invx g1830(.A(n1895), .O(n1894));
  orx  g1831(.A(n1897), .B(n1896), .O(n1895));
  andx g1832(.A(n93), .B(n1900), .O(n1896));
  andx g1833(.A(n1905), .B(n1898), .O(n1897));
  orx  g1834(.A(n1899), .B(n93), .O(n1898));
  andx g1835(.A(n3502), .B(n1900), .O(n1899));
  orx  g1836(.A(n1901), .B(n3480), .O(n1900));
  andx g1837(.A(n3482), .B(n1902), .O(n1901));
  invx g1838(.A(n1903), .O(n1902));
  orx  g1839(.A(n1904), .B(n3521), .O(n1903));
  andx g1840(.A(n1908), .B(pi01), .O(n1904));
  invx g1841(.A(n1906), .O(n1905));
  orx  g1842(.A(n1907), .B(n1912), .O(n1906));
  andx g1843(.A(n1908), .B(n3519), .O(n1907));
  andx g1844(.A(n1909), .B(n93), .O(n1908));
  invx g1845(.A(n1910), .O(n1909));
  andx g1846(.A(n3519), .B(n1911), .O(n1910));
  orx  g1847(.A(n3520), .B(n1912), .O(n1911));
  orx  g1848(.A(n1913), .B(n3495), .O(n1912));
  andx g1849(.A(n1914), .B(n93), .O(n1913));
  andx g1850(.A(pi01), .B(n217), .O(n1914));
  orx  g1851(.A(n1917), .B(n1916), .O(po00));
  andx g1852(.A(n2070), .B(n1919), .O(n1916));
  andx g1853(.A(n1918), .B(n3514), .O(n1917));
  orx  g1854(.A(n2070), .B(n1919), .O(n1918));
  orx  g1855(.A(n1921), .B(n1920), .O(n1919));
  andx g1856(.A(n2063), .B(n1923), .O(n1920));
  andx g1857(.A(n1922), .B(n3529), .O(n1921));
  orx  g1858(.A(n2063), .B(n1923), .O(n1922));
  orx  g1859(.A(n1925), .B(n1924), .O(n1923));
  andx g1860(.A(n2056), .B(n1927), .O(n1924));
  andx g1861(.A(n1926), .B(n141), .O(n1925));
  orx  g1862(.A(n2056), .B(n1927), .O(n1926));
  orx  g1863(.A(n1929), .B(n1928), .O(n1927));
  andx g1864(.A(n2049), .B(n1931), .O(n1928));
  andx g1865(.A(n1930), .B(n144), .O(n1929));
  orx  g1866(.A(n2049), .B(n1931), .O(n1930));
  orx  g1867(.A(n1933), .B(n1932), .O(n1931));
  andx g1868(.A(n2042), .B(n1935), .O(n1932));
  andx g1869(.A(n1934), .B(n198), .O(n1933));
  orx  g1870(.A(n2042), .B(n1935), .O(n1934));
  orx  g1871(.A(n1937), .B(n1936), .O(n1935));
  andx g1872(.A(n2035), .B(n1939), .O(n1936));
  andx g1873(.A(n1938), .B(n208), .O(n1937));
  orx  g1874(.A(n2035), .B(n1939), .O(n1938));
  orx  g1875(.A(n1941), .B(n1940), .O(n1939));
  andx g1876(.A(n2028), .B(n1943), .O(n1940));
  andx g1877(.A(n1942), .B(n213), .O(n1941));
  orx  g1878(.A(n2028), .B(n1943), .O(n1942));
  orx  g1879(.A(n1945), .B(n1944), .O(n1943));
  andx g1880(.A(n2021), .B(n1947), .O(n1944));
  andx g1881(.A(n1946), .B(n113), .O(n1945));
  orx  g1882(.A(n2021), .B(n1947), .O(n1946));
  orx  g1883(.A(n1949), .B(n1948), .O(n1947));
  andx g1884(.A(n2014), .B(n1951), .O(n1948));
  andx g1885(.A(n1950), .B(n118), .O(n1949));
  orx  g1886(.A(n2014), .B(n1951), .O(n1950));
  orx  g1887(.A(n1953), .B(n1952), .O(n1951));
  andx g1888(.A(n2007), .B(n1955), .O(n1952));
  andx g1889(.A(n1954), .B(n120), .O(n1953));
  orx  g1890(.A(n2007), .B(n1955), .O(n1954));
  orx  g1891(.A(n1957), .B(n1956), .O(n1955));
  andx g1892(.A(n2000), .B(n1959), .O(n1956));
  andx g1893(.A(n1958), .B(n95), .O(n1957));
  orx  g1894(.A(n2000), .B(n1959), .O(n1958));
  orx  g1895(.A(n1960), .B(n1961), .O(n1959));
  andx g1896(.A(n1993), .B(n1963), .O(n1960));
  andx g1897(.A(n1962), .B(n130), .O(n1961));
  orx  g1898(.A(n1993), .B(n1963), .O(n1962));
  orx  g1899(.A(n1964), .B(n1965), .O(n1963));
  andx g1900(.A(n1986), .B(n1967), .O(n1964));
  andx g1901(.A(n1966), .B(n103), .O(n1965));
  orx  g1902(.A(n1986), .B(n1967), .O(n1966));
  orx  g1903(.A(n1968), .B(n1969), .O(n1967));
  andx g1904(.A(n1980), .B(n1971), .O(n1968));
  andx g1905(.A(n1970), .B(n105), .O(n1969));
  orx  g1906(.A(n1980), .B(n1971), .O(n1970));
  orx  g1907(.A(n1973), .B(n1972), .O(n1971));
  andx g1908(.A(n1975), .B(n75), .O(n1972));
  andx g1909(.A(n1974), .B(n164), .O(n1973));
  orx  g1910(.A(n75), .B(n1975), .O(n1974));
  orx  g1911(.A(n1977), .B(n1976), .O(n1975));
  andx g1912(.A(n66), .B(n203), .O(n1976));
  andx g1913(.A(pi02), .B(n1978), .O(n1977));
  orx  g1914(.A(n169), .B(n123), .O(n1978));
  orx  g1915(.A(pi00), .B(n123), .O(n1979));
  orx  g1916(.A(n1985), .B(n1981), .O(n1980));
  andx g1917(.A(n1982), .B(n204), .O(n1981));
  andx g1918(.A(n1984), .B(n1983), .O(n1982));
  orx  g1919(.A(n67), .B(n2107), .O(n1983));
  orx  g1920(.A(n66), .B(n2108), .O(n1984));
  andx g1921(.A(n2112), .B(n170), .O(n1985));
  orx  g1922(.A(n1988), .B(n1987), .O(n1986));
  andx g1923(.A(n2121), .B(n169), .O(n1987));
  andx g1924(.A(n1989), .B(n2074), .O(n1988));
  orx  g1925(.A(n1991), .B(n1990), .O(n1989));
  andx g1926(.A(n2117), .B(n2103), .O(n1990));
  andx g1927(.A(n1992), .B(n2116), .O(n1991));
  invx g1928(.A(n2103), .O(n1992));
  orx  g1929(.A(n1995), .B(n1994), .O(n1993));
  andx g1930(.A(n2132), .B(n169), .O(n1994));
  andx g1931(.A(n1996), .B(po02), .O(n1995));
  orx  g1932(.A(n1998), .B(n1997), .O(n1996));
  andx g1933(.A(n2128), .B(n2101), .O(n1997));
  andx g1934(.A(n1999), .B(n2127), .O(n1998));
  invx g1935(.A(n2101), .O(n1999));
  orx  g1936(.A(n2002), .B(n2001), .O(n2000));
  andx g1937(.A(n2144), .B(n170), .O(n2001));
  andx g1938(.A(n2003), .B(n203), .O(n2002));
  orx  g1939(.A(n2005), .B(n2004), .O(n2003));
  andx g1940(.A(n2140), .B(n2099), .O(n2004));
  andx g1941(.A(n2006), .B(n2139), .O(n2005));
  invx g1942(.A(n2099), .O(n2006));
  orx  g1943(.A(n2009), .B(n2008), .O(n2007));
  andx g1944(.A(n2156), .B(n170), .O(n2008));
  andx g1945(.A(n2010), .B(n204), .O(n2009));
  orx  g1946(.A(n2012), .B(n2011), .O(n2010));
  andx g1947(.A(n2152), .B(n2097), .O(n2011));
  andx g1948(.A(n2013), .B(n2151), .O(n2012));
  invx g1949(.A(n2097), .O(n2013));
  orx  g1950(.A(n2016), .B(n2015), .O(n2014));
  andx g1951(.A(n2168), .B(n169), .O(n2015));
  andx g1952(.A(n2017), .B(n204), .O(n2016));
  orx  g1953(.A(n2019), .B(n2018), .O(n2017));
  andx g1954(.A(n2164), .B(n2095), .O(n2018));
  andx g1955(.A(n2020), .B(n2163), .O(n2019));
  invx g1956(.A(n2095), .O(n2020));
  orx  g1957(.A(n2023), .B(n2022), .O(n2021));
  andx g1958(.A(n2180), .B(n170), .O(n2022));
  andx g1959(.A(n2024), .B(po02), .O(n2023));
  orx  g1960(.A(n2026), .B(n2025), .O(n2024));
  andx g1961(.A(n2176), .B(n2093), .O(n2025));
  andx g1962(.A(n2027), .B(n2175), .O(n2026));
  invx g1963(.A(n2093), .O(n2027));
  orx  g1964(.A(n2030), .B(n2029), .O(n2028));
  andx g1965(.A(n2192), .B(n2072), .O(n2029));
  andx g1966(.A(n2031), .B(n203), .O(n2030));
  orx  g1967(.A(n2033), .B(n2032), .O(n2031));
  andx g1968(.A(n2188), .B(n2091), .O(n2032));
  andx g1969(.A(n2034), .B(n2187), .O(n2033));
  invx g1970(.A(n2091), .O(n2034));
  orx  g1971(.A(n2037), .B(n2036), .O(n2035));
  andx g1972(.A(n2204), .B(n169), .O(n2036));
  andx g1973(.A(n2038), .B(n204), .O(n2037));
  orx  g1974(.A(n2040), .B(n2039), .O(n2038));
  andx g1975(.A(n2200), .B(n2089), .O(n2039));
  andx g1976(.A(n2041), .B(n2199), .O(n2040));
  invx g1977(.A(n2089), .O(n2041));
  orx  g1978(.A(n2044), .B(n2043), .O(n2042));
  andx g1979(.A(n2216), .B(n170), .O(n2043));
  andx g1980(.A(n2045), .B(n203), .O(n2044));
  orx  g1981(.A(n2047), .B(n2046), .O(n2045));
  andx g1982(.A(n2212), .B(n2087), .O(n2046));
  andx g1983(.A(n2048), .B(n2211), .O(n2047));
  invx g1984(.A(n2087), .O(n2048));
  orx  g1985(.A(n2051), .B(n2050), .O(n2049));
  andx g1986(.A(n2228), .B(n2072), .O(n2050));
  andx g1987(.A(n2052), .B(po02), .O(n2051));
  orx  g1988(.A(n2054), .B(n2053), .O(n2052));
  andx g1989(.A(n2224), .B(n2085), .O(n2053));
  andx g1990(.A(n2055), .B(n2223), .O(n2054));
  invx g1991(.A(n2085), .O(n2055));
  orx  g1992(.A(n2058), .B(n2057), .O(n2056));
  andx g1993(.A(n2240), .B(n169), .O(n2057));
  andx g1994(.A(n2059), .B(n203), .O(n2058));
  orx  g1995(.A(n2061), .B(n2060), .O(n2059));
  andx g1996(.A(n2236), .B(n2083), .O(n2060));
  andx g1997(.A(n2062), .B(n2235), .O(n2061));
  invx g1998(.A(n2083), .O(n2062));
  orx  g1999(.A(n2065), .B(n2064), .O(n2063));
  andx g2000(.A(n2252), .B(n170), .O(n2064));
  andx g2001(.A(n2066), .B(n204), .O(n2065));
  orx  g2002(.A(n2068), .B(n2067), .O(n2066));
  andx g2003(.A(n2248), .B(n2081), .O(n2067));
  andx g2004(.A(n2069), .B(n2247), .O(n2068));
  invx g2005(.A(n2081), .O(n2069));
  orx  g2006(.A(n2073), .B(n2071), .O(n2070));
  andx g2007(.A(n2264), .B(n2072), .O(n2071));
  invx g2008(.A(po02), .O(n2072));
  andx g2009(.A(n2078), .B(po02), .O(n2073));
  orx  g2010(.A(n2076), .B(n2075), .O(n2074));
  andx g2011(.A(n3513), .B(n2264), .O(n2075));
  andx g2012(.A(n2077), .B(n2260), .O(n2076));
  andx g2013(.A(n2079), .B(n3514), .O(n2077));
  andx g2014(.A(n2259), .B(n2079), .O(n2078));
  orx  g2015(.A(n2080), .B(n2249), .O(n2079));
  andx g2016(.A(n2247), .B(n2081), .O(n2080));
  orx  g2017(.A(n2082), .B(n2237), .O(n2081));
  andx g2018(.A(n2235), .B(n2083), .O(n2082));
  orx  g2019(.A(n2084), .B(n2225), .O(n2083));
  andx g2020(.A(n2223), .B(n2085), .O(n2084));
  orx  g2021(.A(n2086), .B(n2213), .O(n2085));
  andx g2022(.A(n2211), .B(n2087), .O(n2086));
  orx  g2023(.A(n2088), .B(n2201), .O(n2087));
  andx g2024(.A(n2199), .B(n2089), .O(n2088));
  orx  g2025(.A(n2090), .B(n2189), .O(n2089));
  andx g2026(.A(n2187), .B(n2091), .O(n2090));
  orx  g2027(.A(n2092), .B(n2177), .O(n2091));
  andx g2028(.A(n2175), .B(n2093), .O(n2092));
  orx  g2029(.A(n2094), .B(n2165), .O(n2093));
  andx g2030(.A(n2163), .B(n2095), .O(n2094));
  orx  g2031(.A(n2096), .B(n2153), .O(n2095));
  andx g2032(.A(n2151), .B(n2097), .O(n2096));
  orx  g2033(.A(n2098), .B(n2141), .O(n2097));
  andx g2034(.A(n2139), .B(n2099), .O(n2098));
  orx  g2035(.A(n2100), .B(n2129), .O(n2099));
  andx g2036(.A(n2127), .B(n2101), .O(n2100));
  orx  g2037(.A(n2102), .B(n2118), .O(n2101));
  andx g2038(.A(n2116), .B(n2103), .O(n2102));
  orx  g2039(.A(n2105), .B(n2104), .O(n2103));
  andx g2040(.A(n2112), .B(n219), .O(n2104));
  andx g2041(.A(n2107), .B(n67), .O(n2105));
  orx  g2042(.A(pi02), .B(n91), .O(n2106));
  invx g2043(.A(n2108), .O(n2107));
  andx g2044(.A(n2110), .B(n2109), .O(n2108));
  orx  g2045(.A(n2112), .B(pi03), .O(n2109));
  invx g2046(.A(n2111), .O(n2110));
  andx g2047(.A(pi03), .B(n2112), .O(n2111));
  orx  g2048(.A(n2114), .B(n2113), .O(n2112));
  andx g2049(.A(n76), .B(n162), .O(n2113));
  andx g2050(.A(pi04), .B(n2115), .O(n2114));
  orx  g2051(.A(n177), .B(n124), .O(n2115));
  invx g2052(.A(n2117), .O(n2116));
  orx  g2053(.A(n2119), .B(n2118), .O(n2117));
  andx g2054(.A(n2121), .B(n71), .O(n2118));
  invx g2055(.A(n2120), .O(n2119));
  orx  g2056(.A(n2121), .B(n139), .O(n2120));
  orx  g2057(.A(n2126), .B(n2122), .O(n2121));
  andx g2058(.A(n2123), .B(n163), .O(n2122));
  andx g2059(.A(n2125), .B(n2124), .O(n2123));
  orx  g2060(.A(n77), .B(n2299), .O(n2124));
  orx  g2061(.A(n76), .B(n2300), .O(n2125));
  andx g2062(.A(n2304), .B(n178), .O(n2126));
  invx g2063(.A(n2128), .O(n2127));
  orx  g2064(.A(n2130), .B(n2129), .O(n2128));
  andx g2065(.A(n2132), .B(n3517), .O(n2129));
  invx g2066(.A(n2131), .O(n2130));
  orx  g2067(.A(n2132), .B(n134), .O(n2131));
  orx  g2068(.A(n2134), .B(n2133), .O(n2132));
  andx g2069(.A(n2313), .B(n177), .O(n2133));
  andx g2070(.A(n2135), .B(po04), .O(n2134));
  orx  g2071(.A(n2137), .B(n2136), .O(n2135));
  andx g2072(.A(n2309), .B(n2295), .O(n2136));
  andx g2073(.A(n2138), .B(n2308), .O(n2137));
  invx g2074(.A(n2295), .O(n2138));
  invx g2075(.A(n2140), .O(n2139));
  orx  g2076(.A(n2142), .B(n2141), .O(n2140));
  andx g2077(.A(n2144), .B(n130), .O(n2141));
  invx g2078(.A(n2143), .O(n2142));
  orx  g2079(.A(n2144), .B(n3522), .O(n2143));
  orx  g2080(.A(n2146), .B(n2145), .O(n2144));
  andx g2081(.A(n2324), .B(n178), .O(n2145));
  andx g2082(.A(n2147), .B(n162), .O(n2146));
  orx  g2083(.A(n2149), .B(n2148), .O(n2147));
  andx g2084(.A(n2320), .B(n2293), .O(n2148));
  andx g2085(.A(n2150), .B(n2319), .O(n2149));
  invx g2086(.A(n2293), .O(n2150));
  invx g2087(.A(n2152), .O(n2151));
  orx  g2088(.A(n2154), .B(n2153), .O(n2152));
  andx g2089(.A(n2156), .B(n128), .O(n2153));
  invx g2090(.A(n2155), .O(n2154));
  orx  g2091(.A(n73), .B(n2156), .O(n2155));
  orx  g2092(.A(n2158), .B(n2157), .O(n2156));
  andx g2093(.A(n2336), .B(n177), .O(n2157));
  andx g2094(.A(n2159), .B(n163), .O(n2158));
  orx  g2095(.A(n2161), .B(n2160), .O(n2159));
  andx g2096(.A(n2332), .B(n2291), .O(n2160));
  andx g2097(.A(n2162), .B(n2331), .O(n2161));
  invx g2098(.A(n2291), .O(n2162));
  invx g2099(.A(n2164), .O(n2163));
  orx  g2100(.A(n2166), .B(n2165), .O(n2164));
  andx g2101(.A(n2168), .B(n122), .O(n2165));
  invx g2102(.A(n2167), .O(n2166));
  orx  g2103(.A(n122), .B(n2168), .O(n2167));
  orx  g2104(.A(n2170), .B(n2169), .O(n2168));
  andx g2105(.A(n2348), .B(n178), .O(n2169));
  andx g2106(.A(n2171), .B(po04), .O(n2170));
  orx  g2107(.A(n2173), .B(n2172), .O(n2171));
  andx g2108(.A(n2344), .B(n2289), .O(n2172));
  andx g2109(.A(n2174), .B(n2343), .O(n2173));
  invx g2110(.A(n2289), .O(n2174));
  invx g2111(.A(n2176), .O(n2175));
  orx  g2112(.A(n2178), .B(n2177), .O(n2176));
  andx g2113(.A(n2180), .B(n90), .O(n2177));
  invx g2114(.A(n2179), .O(n2178));
  orx  g2115(.A(n117), .B(n2180), .O(n2179));
  orx  g2116(.A(n2182), .B(n2181), .O(n2180));
  andx g2117(.A(n2360), .B(n177), .O(n2181));
  andx g2118(.A(n2183), .B(n162), .O(n2182));
  orx  g2119(.A(n2185), .B(n2184), .O(n2183));
  andx g2120(.A(n2356), .B(n2287), .O(n2184));
  andx g2121(.A(n2186), .B(n2355), .O(n2185));
  invx g2122(.A(n2287), .O(n2186));
  invx g2123(.A(n2188), .O(n2187));
  orx  g2124(.A(n2190), .B(n2189), .O(n2188));
  andx g2125(.A(n2192), .B(n115), .O(n2189));
  invx g2126(.A(n2191), .O(n2190));
  orx  g2127(.A(n3524), .B(n2192), .O(n2191));
  orx  g2128(.A(n2194), .B(n2193), .O(n2192));
  andx g2129(.A(n2372), .B(n178), .O(n2193));
  andx g2130(.A(n2195), .B(n163), .O(n2194));
  orx  g2131(.A(n2197), .B(n2196), .O(n2195));
  andx g2132(.A(n2368), .B(n2285), .O(n2196));
  andx g2133(.A(n2198), .B(n2367), .O(n2197));
  invx g2134(.A(n2285), .O(n2198));
  invx g2135(.A(n2200), .O(n2199));
  orx  g2136(.A(n2202), .B(n2201), .O(n2200));
  andx g2137(.A(n2204), .B(n212), .O(n2201));
  invx g2138(.A(n2203), .O(n2202));
  orx  g2139(.A(n212), .B(n2204), .O(n2203));
  orx  g2140(.A(n2206), .B(n2205), .O(n2204));
  andx g2141(.A(n2384), .B(n177), .O(n2205));
  andx g2142(.A(n2207), .B(po04), .O(n2206));
  orx  g2143(.A(n2209), .B(n2208), .O(n2207));
  andx g2144(.A(n2380), .B(n2283), .O(n2208));
  andx g2145(.A(n2210), .B(n2379), .O(n2209));
  invx g2146(.A(n2283), .O(n2210));
  invx g2147(.A(n2212), .O(n2211));
  orx  g2148(.A(n2214), .B(n2213), .O(n2212));
  andx g2149(.A(n2216), .B(n211), .O(n2213));
  invx g2150(.A(n2215), .O(n2214));
  orx  g2151(.A(n208), .B(n2216), .O(n2215));
  orx  g2152(.A(n2218), .B(n2217), .O(n2216));
  andx g2153(.A(n2396), .B(n178), .O(n2217));
  andx g2154(.A(n2219), .B(n162), .O(n2218));
  orx  g2155(.A(n2221), .B(n2220), .O(n2219));
  andx g2156(.A(n2392), .B(n2281), .O(n2220));
  andx g2157(.A(n2222), .B(n2391), .O(n2221));
  invx g2158(.A(n2281), .O(n2222));
  invx g2159(.A(n2224), .O(n2223));
  orx  g2160(.A(n2226), .B(n2225), .O(n2224));
  andx g2161(.A(n2228), .B(n197), .O(n2225));
  invx g2162(.A(n2227), .O(n2226));
  orx  g2163(.A(n197), .B(n2228), .O(n2227));
  orx  g2164(.A(n2230), .B(n2229), .O(n2228));
  andx g2165(.A(n2408), .B(n177), .O(n2229));
  andx g2166(.A(n2231), .B(n163), .O(n2230));
  orx  g2167(.A(n2233), .B(n2232), .O(n2231));
  andx g2168(.A(n2404), .B(n2279), .O(n2232));
  andx g2169(.A(n2234), .B(n2403), .O(n2233));
  invx g2170(.A(n2279), .O(n2234));
  invx g2171(.A(n2236), .O(n2235));
  orx  g2172(.A(n2238), .B(n2237), .O(n2236));
  andx g2173(.A(n2240), .B(n143), .O(n2237));
  invx g2174(.A(n2239), .O(n2238));
  orx  g2175(.A(n144), .B(n2240), .O(n2239));
  orx  g2176(.A(n2242), .B(n2241), .O(n2240));
  andx g2177(.A(n2420), .B(n178), .O(n2241));
  andx g2178(.A(n2243), .B(po04), .O(n2242));
  orx  g2179(.A(n2245), .B(n2244), .O(n2243));
  andx g2180(.A(n2416), .B(n2277), .O(n2244));
  andx g2181(.A(n2246), .B(n2415), .O(n2245));
  invx g2182(.A(n2277), .O(n2246));
  invx g2183(.A(n2248), .O(n2247));
  orx  g2184(.A(n2250), .B(n2249), .O(n2248));
  andx g2185(.A(n2252), .B(n141), .O(n2249));
  invx g2186(.A(n2251), .O(n2250));
  orx  g2187(.A(n3528), .B(n2252), .O(n2251));
  orx  g2188(.A(n2254), .B(n2253), .O(n2252));
  andx g2189(.A(n2432), .B(n177), .O(n2253));
  andx g2190(.A(n2255), .B(n162), .O(n2254));
  orx  g2191(.A(n2257), .B(n2256), .O(n2255));
  andx g2192(.A(n2428), .B(n2275), .O(n2256));
  andx g2193(.A(n2258), .B(n2427), .O(n2257));
  invx g2194(.A(n2275), .O(n2258));
  invx g2195(.A(n2260), .O(n2259));
  andx g2196(.A(n2263), .B(n2261), .O(n2260));
  invx g2197(.A(n2262), .O(n2261));
  andx g2198(.A(n2264), .B(n3529), .O(n2262));
  orx  g2199(.A(n3529), .B(n2264), .O(n2263));
  orx  g2200(.A(n2267), .B(n2265), .O(n2264));
  andx g2201(.A(n2444), .B(n178), .O(n2265));
  invx g2202(.A(po04), .O(n2266));
  andx g2203(.A(n2272), .B(n163), .O(n2267));
  orx  g2204(.A(n2270), .B(n2269), .O(n2268));
  andx g2205(.A(n3512), .B(n2444), .O(n2269));
  andx g2206(.A(n2271), .B(n2440), .O(n2270));
  andx g2207(.A(n3513), .B(n2273), .O(n2271));
  andx g2208(.A(n2439), .B(n2273), .O(n2272));
  orx  g2209(.A(n2274), .B(n2429), .O(n2273));
  andx g2210(.A(n2427), .B(n2275), .O(n2274));
  orx  g2211(.A(n2276), .B(n2417), .O(n2275));
  andx g2212(.A(n2415), .B(n2277), .O(n2276));
  orx  g2213(.A(n2278), .B(n2405), .O(n2277));
  andx g2214(.A(n2403), .B(n2279), .O(n2278));
  orx  g2215(.A(n2280), .B(n2393), .O(n2279));
  andx g2216(.A(n2391), .B(n2281), .O(n2280));
  orx  g2217(.A(n2282), .B(n2381), .O(n2281));
  andx g2218(.A(n2379), .B(n2283), .O(n2282));
  orx  g2219(.A(n2284), .B(n2369), .O(n2283));
  andx g2220(.A(n2367), .B(n2285), .O(n2284));
  orx  g2221(.A(n2286), .B(n2357), .O(n2285));
  andx g2222(.A(n2355), .B(n2287), .O(n2286));
  orx  g2223(.A(n2288), .B(n2345), .O(n2287));
  andx g2224(.A(n2343), .B(n2289), .O(n2288));
  orx  g2225(.A(n2290), .B(n2333), .O(n2289));
  andx g2226(.A(n2331), .B(n2291), .O(n2290));
  orx  g2227(.A(n2292), .B(n2321), .O(n2291));
  andx g2228(.A(n2319), .B(n2293), .O(n2292));
  orx  g2229(.A(n2294), .B(n2310), .O(n2293));
  andx g2230(.A(n2308), .B(n2295), .O(n2294));
  orx  g2231(.A(n2297), .B(n2296), .O(n2295));
  andx g2232(.A(n2304), .B(n218), .O(n2296));
  andx g2233(.A(n2299), .B(n77), .O(n2297));
  orx  g2234(.A(pi04), .B(n124), .O(n2298));
  invx g2235(.A(n2300), .O(n2299));
  andx g2236(.A(n2302), .B(n2301), .O(n2300));
  orx  g2237(.A(n2304), .B(pi03), .O(n2301));
  invx g2238(.A(n2303), .O(n2302));
  andx g2239(.A(pi03), .B(n2304), .O(n2303));
  orx  g2240(.A(n2306), .B(n2305), .O(n2304));
  andx g2241(.A(n78), .B(n200), .O(n2305));
  andx g2242(.A(pi06), .B(n2307), .O(n2306));
  orx  g2243(.A(n167), .B(n3500), .O(n2307));
  invx g2244(.A(n2309), .O(n2308));
  orx  g2245(.A(n2311), .B(n2310), .O(n2309));
  andx g2246(.A(n2313), .B(n107), .O(n2310));
  invx g2247(.A(n2312), .O(n2311));
  orx  g2248(.A(n2313), .B(n105), .O(n2312));
  orx  g2249(.A(n2318), .B(n2314), .O(n2313));
  andx g2250(.A(n2315), .B(n200), .O(n2314));
  andx g2251(.A(n2317), .B(n2316), .O(n2315));
  orx  g2252(.A(n79), .B(n2477), .O(n2316));
  orx  g2253(.A(n78), .B(n2478), .O(n2317));
  andx g2254(.A(n2482), .B(n167), .O(n2318));
  invx g2255(.A(n2320), .O(n2319));
  orx  g2256(.A(n2322), .B(n2321), .O(n2320));
  andx g2257(.A(n2324), .B(n103), .O(n2321));
  invx g2258(.A(n2323), .O(n2322));
  orx  g2259(.A(n2324), .B(n134), .O(n2323));
  orx  g2260(.A(n2326), .B(n2325), .O(n2324));
  andx g2261(.A(n2491), .B(n168), .O(n2325));
  andx g2262(.A(n2327), .B(n200), .O(n2326));
  orx  g2263(.A(n2329), .B(n2328), .O(n2327));
  andx g2264(.A(n2487), .B(n2473), .O(n2328));
  andx g2265(.A(n2330), .B(n2486), .O(n2329));
  invx g2266(.A(n2473), .O(n2330));
  invx g2267(.A(n2332), .O(n2331));
  orx  g2268(.A(n2334), .B(n2333), .O(n2332));
  andx g2269(.A(n2336), .B(n130), .O(n2333));
  invx g2270(.A(n2335), .O(n2334));
  orx  g2271(.A(n2336), .B(n130), .O(n2335));
  orx  g2272(.A(n2338), .B(n2337), .O(n2336));
  andx g2273(.A(n2502), .B(n167), .O(n2337));
  andx g2274(.A(n2339), .B(n201), .O(n2338));
  orx  g2275(.A(n2341), .B(n2340), .O(n2339));
  andx g2276(.A(n2498), .B(n2471), .O(n2340));
  andx g2277(.A(n2342), .B(n2497), .O(n2341));
  invx g2278(.A(n2471), .O(n2342));
  invx g2279(.A(n2344), .O(n2343));
  orx  g2280(.A(n2346), .B(n2345), .O(n2344));
  andx g2281(.A(n2348), .B(n95), .O(n2345));
  invx g2282(.A(n2347), .O(n2346));
  orx  g2283(.A(n129), .B(n2348), .O(n2347));
  orx  g2284(.A(n2350), .B(n2349), .O(n2348));
  andx g2285(.A(n2514), .B(n168), .O(n2349));
  andx g2286(.A(n2351), .B(po06), .O(n2350));
  orx  g2287(.A(n2353), .B(n2352), .O(n2351));
  andx g2288(.A(n2510), .B(n2469), .O(n2352));
  andx g2289(.A(n2354), .B(n2509), .O(n2353));
  invx g2290(.A(n2469), .O(n2354));
  invx g2291(.A(n2356), .O(n2355));
  orx  g2292(.A(n2358), .B(n2357), .O(n2356));
  andx g2293(.A(n2360), .B(n72), .O(n2357));
  invx g2294(.A(n2359), .O(n2358));
  orx  g2295(.A(n72), .B(n2360), .O(n2359));
  orx  g2296(.A(n2362), .B(n2361), .O(n2360));
  andx g2297(.A(n2526), .B(n167), .O(n2361));
  andx g2298(.A(n2363), .B(n201), .O(n2362));
  orx  g2299(.A(n2365), .B(n2364), .O(n2363));
  andx g2300(.A(n2522), .B(n2467), .O(n2364));
  andx g2301(.A(n2366), .B(n2521), .O(n2365));
  invx g2302(.A(n2467), .O(n2366));
  invx g2303(.A(n2368), .O(n2367));
  orx  g2304(.A(n2370), .B(n2369), .O(n2368));
  andx g2305(.A(n2372), .B(n118), .O(n2369));
  invx g2306(.A(n2371), .O(n2370));
  orx  g2307(.A(n117), .B(n2372), .O(n2371));
  orx  g2308(.A(n2374), .B(n2373), .O(n2372));
  andx g2309(.A(n2538), .B(n168), .O(n2373));
  andx g2310(.A(n2375), .B(po06), .O(n2374));
  orx  g2311(.A(n2377), .B(n2376), .O(n2375));
  andx g2312(.A(n2534), .B(n2465), .O(n2376));
  andx g2313(.A(n2378), .B(n2533), .O(n2377));
  invx g2314(.A(n2465), .O(n2378));
  invx g2315(.A(n2380), .O(n2379));
  orx  g2316(.A(n2382), .B(n2381), .O(n2380));
  andx g2317(.A(n2384), .B(n115), .O(n2381));
  invx g2318(.A(n2383), .O(n2382));
  orx  g2319(.A(n114), .B(n2384), .O(n2383));
  orx  g2320(.A(n2386), .B(n2385), .O(n2384));
  andx g2321(.A(n2550), .B(n167), .O(n2385));
  andx g2322(.A(n2387), .B(n201), .O(n2386));
  orx  g2323(.A(n2389), .B(n2388), .O(n2387));
  andx g2324(.A(n2546), .B(n2463), .O(n2388));
  andx g2325(.A(n2390), .B(n2545), .O(n2389));
  invx g2326(.A(n2463), .O(n2390));
  invx g2327(.A(n2392), .O(n2391));
  orx  g2328(.A(n2394), .B(n2393), .O(n2392));
  andx g2329(.A(n2396), .B(n215), .O(n2393));
  invx g2330(.A(n2395), .O(n2394));
  orx  g2331(.A(n215), .B(n2396), .O(n2395));
  orx  g2332(.A(n2398), .B(n2397), .O(n2396));
  andx g2333(.A(n2562), .B(n168), .O(n2397));
  andx g2334(.A(n2399), .B(n200), .O(n2398));
  orx  g2335(.A(n2401), .B(n2400), .O(n2399));
  andx g2336(.A(n2558), .B(n2461), .O(n2400));
  andx g2337(.A(n2402), .B(n2557), .O(n2401));
  invx g2338(.A(n2461), .O(n2402));
  invx g2339(.A(n2404), .O(n2403));
  orx  g2340(.A(n2406), .B(n2405), .O(n2404));
  andx g2341(.A(n2408), .B(n210), .O(n2405));
  invx g2342(.A(n2407), .O(n2406));
  orx  g2343(.A(n211), .B(n2408), .O(n2407));
  orx  g2344(.A(n2410), .B(n2409), .O(n2408));
  andx g2345(.A(n2574), .B(n167), .O(n2409));
  andx g2346(.A(n2411), .B(n201), .O(n2410));
  orx  g2347(.A(n2413), .B(n2412), .O(n2411));
  andx g2348(.A(n2570), .B(n2459), .O(n2412));
  andx g2349(.A(n2414), .B(n2569), .O(n2413));
  invx g2350(.A(n2459), .O(n2414));
  invx g2351(.A(n2416), .O(n2415));
  orx  g2352(.A(n2418), .B(n2417), .O(n2416));
  andx g2353(.A(n2420), .B(n199), .O(n2417));
  invx g2354(.A(n2419), .O(n2418));
  orx  g2355(.A(n199), .B(n2420), .O(n2419));
  orx  g2356(.A(n2422), .B(n2421), .O(n2420));
  andx g2357(.A(n2586), .B(n168), .O(n2421));
  andx g2358(.A(n2423), .B(n201), .O(n2422));
  orx  g2359(.A(n2425), .B(n2424), .O(n2423));
  andx g2360(.A(n2582), .B(n2457), .O(n2424));
  andx g2361(.A(n2426), .B(n2581), .O(n2425));
  invx g2362(.A(n2457), .O(n2426));
  invx g2363(.A(n2428), .O(n2427));
  orx  g2364(.A(n2430), .B(n2429), .O(n2428));
  andx g2365(.A(n2432), .B(n144), .O(n2429));
  invx g2366(.A(n2431), .O(n2430));
  orx  g2367(.A(n3527), .B(n2432), .O(n2431));
  orx  g2368(.A(n2434), .B(n2433), .O(n2432));
  andx g2369(.A(n2598), .B(n167), .O(n2433));
  andx g2370(.A(n2435), .B(n201), .O(n2434));
  orx  g2371(.A(n2437), .B(n2436), .O(n2435));
  andx g2372(.A(n2594), .B(n2455), .O(n2436));
  andx g2373(.A(n2438), .B(n2593), .O(n2437));
  invx g2374(.A(n2455), .O(n2438));
  invx g2375(.A(n2440), .O(n2439));
  andx g2376(.A(n2443), .B(n2441), .O(n2440));
  invx g2377(.A(n2442), .O(n2441));
  andx g2378(.A(n2444), .B(n3528), .O(n2442));
  orx  g2379(.A(n3528), .B(n2444), .O(n2443));
  orx  g2380(.A(n2447), .B(n2445), .O(n2444));
  andx g2381(.A(n2610), .B(n168), .O(n2445));
  invx g2382(.A(n200), .O(n2446));
  andx g2383(.A(n2452), .B(n200), .O(n2447));
  orx  g2384(.A(n2450), .B(n2449), .O(po06));
  andx g2385(.A(n3511), .B(n2610), .O(n2449));
  andx g2386(.A(n2451), .B(n2606), .O(n2450));
  andx g2387(.A(n3512), .B(n2453), .O(n2451));
  andx g2388(.A(n2605), .B(n2453), .O(n2452));
  orx  g2389(.A(n2454), .B(n2595), .O(n2453));
  andx g2390(.A(n2593), .B(n2455), .O(n2454));
  orx  g2391(.A(n2456), .B(n2583), .O(n2455));
  andx g2392(.A(n2581), .B(n2457), .O(n2456));
  orx  g2393(.A(n2458), .B(n2571), .O(n2457));
  andx g2394(.A(n2569), .B(n2459), .O(n2458));
  orx  g2395(.A(n2460), .B(n2559), .O(n2459));
  andx g2396(.A(n2557), .B(n2461), .O(n2460));
  orx  g2397(.A(n2462), .B(n2547), .O(n2461));
  andx g2398(.A(n2545), .B(n2463), .O(n2462));
  orx  g2399(.A(n2464), .B(n2535), .O(n2463));
  andx g2400(.A(n2533), .B(n2465), .O(n2464));
  orx  g2401(.A(n2466), .B(n2523), .O(n2465));
  andx g2402(.A(n2521), .B(n2467), .O(n2466));
  orx  g2403(.A(n2468), .B(n2511), .O(n2467));
  andx g2404(.A(n2509), .B(n2469), .O(n2468));
  orx  g2405(.A(n2470), .B(n2499), .O(n2469));
  andx g2406(.A(n2497), .B(n2471), .O(n2470));
  orx  g2407(.A(n2472), .B(n2488), .O(n2471));
  andx g2408(.A(n2486), .B(n2473), .O(n2472));
  orx  g2409(.A(n2475), .B(n2474), .O(n2473));
  andx g2410(.A(n2482), .B(n216), .O(n2474));
  andx g2411(.A(n2477), .B(n79), .O(n2475));
  orx  g2412(.A(pi06), .B(n126), .O(n2476));
  invx g2413(.A(n2478), .O(n2477));
  andx g2414(.A(n2480), .B(n2479), .O(n2478));
  orx  g2415(.A(n2482), .B(pi03), .O(n2479));
  invx g2416(.A(n2481), .O(n2480));
  andx g2417(.A(pi03), .B(n2482), .O(n2481));
  orx  g2418(.A(n2484), .B(n2483), .O(n2482));
  andx g2419(.A(n68), .B(n159), .O(n2483));
  andx g2420(.A(pi08), .B(n2485), .O(n2484));
  orx  g2421(.A(n2612), .B(n126), .O(n2485));
  invx g2422(.A(n2487), .O(n2486));
  orx  g2423(.A(n2489), .B(n2488), .O(n2487));
  andx g2424(.A(n2491), .B(n105), .O(n2488));
  invx g2425(.A(n2490), .O(n2489));
  orx  g2426(.A(n2491), .B(n108), .O(n2490));
  orx  g2427(.A(n2496), .B(n2492), .O(n2491));
  andx g2428(.A(n2493), .B(n159), .O(n2492));
  andx g2429(.A(n2495), .B(n2494), .O(n2493));
  orx  g2430(.A(n69), .B(n2641), .O(n2494));
  orx  g2431(.A(n68), .B(n2642), .O(n2495));
  andx g2432(.A(n2646), .B(n148), .O(n2496));
  invx g2433(.A(n2498), .O(n2497));
  orx  g2434(.A(n2500), .B(n2499), .O(n2498));
  andx g2435(.A(n2502), .B(n103), .O(n2499));
  invx g2436(.A(n2501), .O(n2500));
  orx  g2437(.A(n2502), .B(n135), .O(n2501));
  orx  g2438(.A(n2504), .B(n2503), .O(n2502));
  andx g2439(.A(n2655), .B(n148), .O(n2503));
  andx g2440(.A(n2505), .B(n159), .O(n2504));
  orx  g2441(.A(n2507), .B(n2506), .O(n2505));
  andx g2442(.A(n2651), .B(n2637), .O(n2506));
  andx g2443(.A(n2508), .B(n2650), .O(n2507));
  invx g2444(.A(n2637), .O(n2508));
  invx g2445(.A(n2510), .O(n2509));
  orx  g2446(.A(n2512), .B(n2511), .O(n2510));
  andx g2447(.A(n2514), .B(n131), .O(n2511));
  invx g2448(.A(n2513), .O(n2512));
  orx  g2449(.A(n2514), .B(n130), .O(n2513));
  orx  g2450(.A(n2516), .B(n2515), .O(n2514));
  andx g2451(.A(n2666), .B(n148), .O(n2515));
  andx g2452(.A(n2517), .B(po08), .O(n2516));
  orx  g2453(.A(n2519), .B(n2518), .O(n2517));
  andx g2454(.A(n2662), .B(n2635), .O(n2518));
  andx g2455(.A(n2520), .B(n2661), .O(n2519));
  invx g2456(.A(n2635), .O(n2520));
  invx g2457(.A(n2522), .O(n2521));
  orx  g2458(.A(n2524), .B(n2523), .O(n2522));
  andx g2459(.A(n2526), .B(n128), .O(n2523));
  invx g2460(.A(n2525), .O(n2524));
  orx  g2461(.A(n96), .B(n2526), .O(n2525));
  orx  g2462(.A(n2528), .B(n2527), .O(n2526));
  andx g2463(.A(n2678), .B(n148), .O(n2527));
  andx g2464(.A(n2529), .B(n2614), .O(n2528));
  orx  g2465(.A(n2531), .B(n2530), .O(n2529));
  andx g2466(.A(n2674), .B(n2633), .O(n2530));
  andx g2467(.A(n2532), .B(n2673), .O(n2531));
  invx g2468(.A(n2633), .O(n2532));
  invx g2469(.A(n2534), .O(n2533));
  orx  g2470(.A(n2536), .B(n2535), .O(n2534));
  andx g2471(.A(n2538), .B(n122), .O(n2535));
  invx g2472(.A(n2537), .O(n2536));
  orx  g2473(.A(n120), .B(n2538), .O(n2537));
  orx  g2474(.A(n2540), .B(n2539), .O(n2538));
  andx g2475(.A(n2690), .B(n148), .O(n2539));
  andx g2476(.A(n2541), .B(po08), .O(n2540));
  orx  g2477(.A(n2543), .B(n2542), .O(n2541));
  andx g2478(.A(n2686), .B(n2631), .O(n2542));
  andx g2479(.A(n2544), .B(n2685), .O(n2543));
  invx g2480(.A(n2631), .O(n2544));
  invx g2481(.A(n2546), .O(n2545));
  orx  g2482(.A(n2548), .B(n2547), .O(n2546));
  andx g2483(.A(n2550), .B(n117), .O(n2547));
  invx g2484(.A(n2549), .O(n2548));
  orx  g2485(.A(n117), .B(n2550), .O(n2549));
  orx  g2486(.A(n2552), .B(n2551), .O(n2550));
  andx g2487(.A(n2702), .B(n148), .O(n2551));
  andx g2488(.A(n2553), .B(n2614), .O(n2552));
  orx  g2489(.A(n2555), .B(n2554), .O(n2553));
  andx g2490(.A(n2698), .B(n2629), .O(n2554));
  andx g2491(.A(n2556), .B(n2697), .O(n2555));
  invx g2492(.A(n2629), .O(n2556));
  invx g2493(.A(n2558), .O(n2557));
  orx  g2494(.A(n2560), .B(n2559), .O(n2558));
  andx g2495(.A(n2562), .B(n115), .O(n2559));
  invx g2496(.A(n2561), .O(n2560));
  orx  g2497(.A(n114), .B(n2562), .O(n2561));
  orx  g2498(.A(n2564), .B(n2563), .O(n2562));
  andx g2499(.A(n2714), .B(n2612), .O(n2563));
  andx g2500(.A(n2565), .B(po08), .O(n2564));
  orx  g2501(.A(n2567), .B(n2566), .O(n2565));
  andx g2502(.A(n2710), .B(n2627), .O(n2566));
  andx g2503(.A(n2568), .B(n2709), .O(n2567));
  invx g2504(.A(n2627), .O(n2568));
  invx g2505(.A(n2570), .O(n2569));
  orx  g2506(.A(n2572), .B(n2571), .O(n2570));
  andx g2507(.A(n2574), .B(n214), .O(n2571));
  invx g2508(.A(n2573), .O(n2572));
  orx  g2509(.A(n214), .B(n2574), .O(n2573));
  orx  g2510(.A(n2576), .B(n2575), .O(n2574));
  andx g2511(.A(n2726), .B(n2612), .O(n2575));
  andx g2512(.A(n2577), .B(n159), .O(n2576));
  orx  g2513(.A(n2579), .B(n2578), .O(n2577));
  andx g2514(.A(n2722), .B(n2625), .O(n2578));
  andx g2515(.A(n2580), .B(n2721), .O(n2579));
  invx g2516(.A(n2625), .O(n2580));
  invx g2517(.A(n2582), .O(n2581));
  orx  g2518(.A(n2584), .B(n2583), .O(n2582));
  andx g2519(.A(n2586), .B(n209), .O(n2583));
  invx g2520(.A(n2585), .O(n2584));
  orx  g2521(.A(n210), .B(n2586), .O(n2585));
  orx  g2522(.A(n2588), .B(n2587), .O(n2586));
  andx g2523(.A(n2738), .B(n2612), .O(n2587));
  andx g2524(.A(n2589), .B(po08), .O(n2588));
  orx  g2525(.A(n2591), .B(n2590), .O(n2589));
  andx g2526(.A(n2734), .B(n2623), .O(n2590));
  andx g2527(.A(n2592), .B(n2733), .O(n2591));
  invx g2528(.A(n2623), .O(n2592));
  invx g2529(.A(n2594), .O(n2593));
  orx  g2530(.A(n2596), .B(n2595), .O(n2594));
  andx g2531(.A(n2598), .B(n198), .O(n2595));
  invx g2532(.A(n2597), .O(n2596));
  orx  g2533(.A(n198), .B(n2598), .O(n2597));
  orx  g2534(.A(n2600), .B(n2599), .O(n2598));
  andx g2535(.A(n2750), .B(n2612), .O(n2599));
  andx g2536(.A(n2601), .B(po08), .O(n2600));
  orx  g2537(.A(n2603), .B(n2602), .O(n2601));
  andx g2538(.A(n2746), .B(n2621), .O(n2602));
  andx g2539(.A(n2604), .B(n2745), .O(n2603));
  invx g2540(.A(n2621), .O(n2604));
  invx g2541(.A(n2606), .O(n2605));
  andx g2542(.A(n2609), .B(n2607), .O(n2606));
  invx g2543(.A(n2608), .O(n2607));
  andx g2544(.A(n2610), .B(n3527), .O(n2608));
  orx  g2545(.A(n143), .B(n2610), .O(n2609));
  orx  g2546(.A(n2613), .B(n2611), .O(n2610));
  andx g2547(.A(n2762), .B(n2612), .O(n2611));
  invx g2548(.A(n159), .O(n2612));
  andx g2549(.A(n2618), .B(po08), .O(n2613));
  orx  g2550(.A(n2616), .B(n2615), .O(n2614));
  andx g2551(.A(n3510), .B(n2762), .O(n2615));
  andx g2552(.A(n2617), .B(n2758), .O(n2616));
  andx g2553(.A(n3511), .B(n2619), .O(n2617));
  andx g2554(.A(n2757), .B(n2619), .O(n2618));
  orx  g2555(.A(n2620), .B(n2747), .O(n2619));
  andx g2556(.A(n2745), .B(n2621), .O(n2620));
  orx  g2557(.A(n2622), .B(n2735), .O(n2621));
  andx g2558(.A(n2733), .B(n2623), .O(n2622));
  orx  g2559(.A(n2624), .B(n2723), .O(n2623));
  andx g2560(.A(n2721), .B(n2625), .O(n2624));
  orx  g2561(.A(n2626), .B(n2711), .O(n2625));
  andx g2562(.A(n2709), .B(n2627), .O(n2626));
  orx  g2563(.A(n2628), .B(n2699), .O(n2627));
  andx g2564(.A(n2697), .B(n2629), .O(n2628));
  orx  g2565(.A(n2630), .B(n2687), .O(n2629));
  andx g2566(.A(n2685), .B(n2631), .O(n2630));
  orx  g2567(.A(n2632), .B(n2675), .O(n2631));
  andx g2568(.A(n2673), .B(n2633), .O(n2632));
  orx  g2569(.A(n2634), .B(n2663), .O(n2633));
  andx g2570(.A(n2661), .B(n2635), .O(n2634));
  orx  g2571(.A(n2636), .B(n2652), .O(n2635));
  andx g2572(.A(n2650), .B(n2637), .O(n2636));
  orx  g2573(.A(n2639), .B(n2638), .O(n2637));
  andx g2574(.A(n2646), .B(n164), .O(n2638));
  andx g2575(.A(n2641), .B(n69), .O(n2639));
  orx  g2576(.A(pi08), .B(n3500), .O(n2640));
  invx g2577(.A(n2642), .O(n2641));
  andx g2578(.A(n2644), .B(n2643), .O(n2642));
  orx  g2579(.A(n2646), .B(pi03), .O(n2643));
  invx g2580(.A(n2645), .O(n2644));
  andx g2581(.A(pi03), .B(n2646), .O(n2645));
  orx  g2582(.A(n2648), .B(n2647), .O(n2646));
  andx g2583(.A(n88), .B(n180), .O(n2647));
  andx g2584(.A(pi10), .B(n2649), .O(n2648));
  orx  g2585(.A(n2764), .B(n125), .O(n2649));
  invx g2586(.A(n2651), .O(n2650));
  orx  g2587(.A(n2653), .B(n2652), .O(n2651));
  andx g2588(.A(n2655), .B(n139), .O(n2652));
  invx g2589(.A(n2654), .O(n2653));
  orx  g2590(.A(n2655), .B(n3518), .O(n2654));
  orx  g2591(.A(n2660), .B(n2656), .O(n2655));
  andx g2592(.A(n2657), .B(n2766), .O(n2656));
  andx g2593(.A(n2659), .B(n2658), .O(n2657));
  orx  g2594(.A(n89), .B(n2791), .O(n2658));
  orx  g2595(.A(n88), .B(n2792), .O(n2659));
  andx g2596(.A(n2796), .B(n147), .O(n2660));
  invx g2597(.A(n2662), .O(n2661));
  orx  g2598(.A(n2664), .B(n2663), .O(n2662));
  andx g2599(.A(n2666), .B(n133), .O(n2663));
  invx g2600(.A(n2665), .O(n2664));
  orx  g2601(.A(n2666), .B(n103), .O(n2665));
  orx  g2602(.A(n2668), .B(n2667), .O(n2666));
  andx g2603(.A(n2805), .B(n147), .O(n2667));
  andx g2604(.A(n2669), .B(po10), .O(n2668));
  orx  g2605(.A(n2671), .B(n2670), .O(n2669));
  andx g2606(.A(n2801), .B(n2787), .O(n2670));
  andx g2607(.A(n2672), .B(n2800), .O(n2671));
  invx g2608(.A(n2787), .O(n2672));
  invx g2609(.A(n2674), .O(n2673));
  orx  g2610(.A(n2676), .B(n2675), .O(n2674));
  andx g2611(.A(n2678), .B(n131), .O(n2675));
  invx g2612(.A(n2677), .O(n2676));
  orx  g2613(.A(n2678), .B(n130), .O(n2677));
  orx  g2614(.A(n2680), .B(n2679), .O(n2678));
  andx g2615(.A(n2816), .B(n147), .O(n2679));
  andx g2616(.A(n2681), .B(n180), .O(n2680));
  orx  g2617(.A(n2683), .B(n2682), .O(n2681));
  andx g2618(.A(n2812), .B(n2785), .O(n2682));
  andx g2619(.A(n2684), .B(n2811), .O(n2683));
  invx g2620(.A(n2785), .O(n2684));
  invx g2621(.A(n2686), .O(n2685));
  orx  g2622(.A(n2688), .B(n2687), .O(n2686));
  andx g2623(.A(n2690), .B(n129), .O(n2687));
  invx g2624(.A(n2689), .O(n2688));
  orx  g2625(.A(n129), .B(n2690), .O(n2689));
  orx  g2626(.A(n2692), .B(n2691), .O(n2690));
  andx g2627(.A(n2828), .B(n147), .O(n2691));
  andx g2628(.A(n2693), .B(n2766), .O(n2692));
  orx  g2629(.A(n2695), .B(n2694), .O(n2693));
  andx g2630(.A(n2824), .B(n2783), .O(n2694));
  andx g2631(.A(n2696), .B(n2823), .O(n2695));
  invx g2632(.A(n2783), .O(n2696));
  invx g2633(.A(n2698), .O(n2697));
  orx  g2634(.A(n2700), .B(n2699), .O(n2698));
  andx g2635(.A(n2702), .B(n72), .O(n2699));
  invx g2636(.A(n2701), .O(n2700));
  orx  g2637(.A(n122), .B(n2702), .O(n2701));
  orx  g2638(.A(n2704), .B(n2703), .O(n2702));
  andx g2639(.A(n2840), .B(n147), .O(n2703));
  andx g2640(.A(n2705), .B(po10), .O(n2704));
  orx  g2641(.A(n2707), .B(n2706), .O(n2705));
  andx g2642(.A(n2836), .B(n2781), .O(n2706));
  andx g2643(.A(n2708), .B(n2835), .O(n2707));
  invx g2644(.A(n2781), .O(n2708));
  invx g2645(.A(n2710), .O(n2709));
  orx  g2646(.A(n2712), .B(n2711), .O(n2710));
  andx g2647(.A(n2714), .B(n116), .O(n2711));
  invx g2648(.A(n2713), .O(n2712));
  orx  g2649(.A(n3523), .B(n2714), .O(n2713));
  orx  g2650(.A(n2716), .B(n2715), .O(n2714));
  andx g2651(.A(n2852), .B(n2764), .O(n2715));
  andx g2652(.A(n2717), .B(n180), .O(n2716));
  orx  g2653(.A(n2719), .B(n2718), .O(n2717));
  andx g2654(.A(n2848), .B(n2779), .O(n2718));
  andx g2655(.A(n2720), .B(n2847), .O(n2719));
  invx g2656(.A(n2779), .O(n2720));
  invx g2657(.A(n2722), .O(n2721));
  orx  g2658(.A(n2724), .B(n2723), .O(n2722));
  andx g2659(.A(n2726), .B(n3524), .O(n2723));
  invx g2660(.A(n2725), .O(n2724));
  orx  g2661(.A(n115), .B(n2726), .O(n2725));
  orx  g2662(.A(n2728), .B(n2727), .O(n2726));
  andx g2663(.A(n2864), .B(n2764), .O(n2727));
  andx g2664(.A(n2729), .B(n180), .O(n2728));
  orx  g2665(.A(n2731), .B(n2730), .O(n2729));
  andx g2666(.A(n2860), .B(n2777), .O(n2730));
  andx g2667(.A(n2732), .B(n2859), .O(n2731));
  invx g2668(.A(n2777), .O(n2732));
  invx g2669(.A(n2734), .O(n2733));
  orx  g2670(.A(n2736), .B(n2735), .O(n2734));
  andx g2671(.A(n2738), .B(n213), .O(n2735));
  invx g2672(.A(n2737), .O(n2736));
  orx  g2673(.A(n213), .B(n2738), .O(n2737));
  orx  g2674(.A(n2740), .B(n2739), .O(n2738));
  andx g2675(.A(n2876), .B(n2764), .O(n2739));
  andx g2676(.A(n2741), .B(po10), .O(n2740));
  orx  g2677(.A(n2743), .B(n2742), .O(n2741));
  andx g2678(.A(n2872), .B(n2775), .O(n2742));
  andx g2679(.A(n2744), .B(n2871), .O(n2743));
  invx g2680(.A(n2775), .O(n2744));
  invx g2681(.A(n2746), .O(n2745));
  orx  g2682(.A(n2748), .B(n2747), .O(n2746));
  andx g2683(.A(n2750), .B(n208), .O(n2747));
  invx g2684(.A(n2749), .O(n2748));
  orx  g2685(.A(n209), .B(n2750), .O(n2749));
  orx  g2686(.A(n2752), .B(n2751), .O(n2750));
  andx g2687(.A(n2888), .B(n2764), .O(n2751));
  andx g2688(.A(n2753), .B(n180), .O(n2752));
  orx  g2689(.A(n2755), .B(n2754), .O(n2753));
  andx g2690(.A(n2884), .B(n2773), .O(n2754));
  andx g2691(.A(n2756), .B(n2883), .O(n2755));
  invx g2692(.A(n2773), .O(n2756));
  invx g2693(.A(n2758), .O(n2757));
  andx g2694(.A(n2761), .B(n2759), .O(n2758));
  invx g2695(.A(n2760), .O(n2759));
  andx g2696(.A(n2762), .B(n197), .O(n2760));
  orx  g2697(.A(n197), .B(n2762), .O(n2761));
  orx  g2698(.A(n2765), .B(n2763), .O(n2762));
  andx g2699(.A(n2900), .B(n2764), .O(n2763));
  invx g2700(.A(po10), .O(n2764));
  andx g2701(.A(n2770), .B(po10), .O(n2765));
  orx  g2702(.A(n2768), .B(n2767), .O(n2766));
  andx g2703(.A(n3509), .B(n2900), .O(n2767));
  andx g2704(.A(n2769), .B(n2896), .O(n2768));
  andx g2705(.A(n3510), .B(n2771), .O(n2769));
  andx g2706(.A(n2895), .B(n2771), .O(n2770));
  orx  g2707(.A(n2772), .B(n2885), .O(n2771));
  andx g2708(.A(n2883), .B(n2773), .O(n2772));
  orx  g2709(.A(n2774), .B(n2873), .O(n2773));
  andx g2710(.A(n2871), .B(n2775), .O(n2774));
  orx  g2711(.A(n2776), .B(n2861), .O(n2775));
  andx g2712(.A(n2859), .B(n2777), .O(n2776));
  orx  g2713(.A(n2778), .B(n2849), .O(n2777));
  andx g2714(.A(n2847), .B(n2779), .O(n2778));
  orx  g2715(.A(n2780), .B(n2837), .O(n2779));
  andx g2716(.A(n2835), .B(n2781), .O(n2780));
  orx  g2717(.A(n2782), .B(n2825), .O(n2781));
  andx g2718(.A(n2823), .B(n2783), .O(n2782));
  orx  g2719(.A(n2784), .B(n2813), .O(n2783));
  andx g2720(.A(n2811), .B(n2785), .O(n2784));
  orx  g2721(.A(n2786), .B(n2802), .O(n2785));
  andx g2722(.A(n2800), .B(n2787), .O(n2786));
  orx  g2723(.A(n2789), .B(n2788), .O(n2787));
  andx g2724(.A(n2796), .B(n219), .O(n2788));
  andx g2725(.A(n2791), .B(n89), .O(n2789));
  orx  g2726(.A(pi10), .B(n125), .O(n2790));
  invx g2727(.A(n2792), .O(n2791));
  andx g2728(.A(n2794), .B(n2793), .O(n2792));
  orx  g2729(.A(n2796), .B(pi03), .O(n2793));
  invx g2730(.A(n2795), .O(n2794));
  andx g2731(.A(pi03), .B(n2796), .O(n2795));
  orx  g2732(.A(n2798), .B(n2797), .O(n2796));
  andx g2733(.A(po12), .B(n64), .O(n2797));
  andx g2734(.A(pi12), .B(n2799), .O(n2798));
  orx  g2735(.A(n125), .B(n157), .O(n2799));
  invx g2736(.A(n2801), .O(n2800));
  orx  g2737(.A(n2803), .B(n2802), .O(n2801));
  andx g2738(.A(n2805), .B(n105), .O(n2802));
  invx g2739(.A(n2804), .O(n2803));
  orx  g2740(.A(n2805), .B(n137), .O(n2804));
  orx  g2741(.A(n2810), .B(n2806), .O(n2805));
  andx g2742(.A(n2807), .B(po12), .O(n2806));
  andx g2743(.A(n2809), .B(n2808), .O(n2807));
  orx  g2744(.A(n65), .B(n2931), .O(n2808));
  orx  g2745(.A(n64), .B(n2932), .O(n2809));
  andx g2746(.A(n2936), .B(n158), .O(n2810));
  invx g2747(.A(n2812), .O(n2811));
  orx  g2748(.A(n2814), .B(n2813), .O(n2812));
  andx g2749(.A(n2816), .B(n104), .O(n2813));
  invx g2750(.A(n2815), .O(n2814));
  orx  g2751(.A(n2816), .B(n3517), .O(n2815));
  orx  g2752(.A(n2822), .B(n2817), .O(n2816));
  andx g2753(.A(n2818), .B(n2902), .O(n2817));
  orx  g2754(.A(n2820), .B(n2819), .O(n2818));
  andx g2755(.A(n2941), .B(n2927), .O(n2819));
  andx g2756(.A(n2821), .B(n2940), .O(n2820));
  invx g2757(.A(n2927), .O(n2821));
  andx g2758(.A(n2945), .B(n157), .O(n2822));
  invx g2759(.A(n2824), .O(n2823));
  orx  g2760(.A(n2826), .B(n2825), .O(n2824));
  andx g2761(.A(n2828), .B(n131), .O(n2825));
  invx g2762(.A(n2827), .O(n2826));
  orx  g2763(.A(n2828), .B(n3522), .O(n2827));
  orx  g2764(.A(n2834), .B(n2829), .O(n2828));
  andx g2765(.A(n2830), .B(po12), .O(n2829));
  orx  g2766(.A(n2832), .B(n2831), .O(n2830));
  andx g2767(.A(n2952), .B(n2925), .O(n2831));
  andx g2768(.A(n2833), .B(n2951), .O(n2832));
  invx g2769(.A(n2925), .O(n2833));
  andx g2770(.A(n2956), .B(n158), .O(n2834));
  invx g2771(.A(n2836), .O(n2835));
  orx  g2772(.A(n2838), .B(n2837), .O(n2836));
  andx g2773(.A(n2840), .B(n73), .O(n2837));
  invx g2774(.A(n2839), .O(n2838));
  orx  g2775(.A(n127), .B(n2840), .O(n2839));
  orx  g2776(.A(n2846), .B(n2841), .O(n2840));
  andx g2777(.A(n2842), .B(n2902), .O(n2841));
  orx  g2778(.A(n2844), .B(n2843), .O(n2842));
  andx g2779(.A(n2964), .B(n2923), .O(n2843));
  andx g2780(.A(n2845), .B(n2963), .O(n2844));
  invx g2781(.A(n2923), .O(n2845));
  andx g2782(.A(n2968), .B(n157), .O(n2846));
  invx g2783(.A(n2848), .O(n2847));
  orx  g2784(.A(n2850), .B(n2849), .O(n2848));
  andx g2785(.A(n2852), .B(n94), .O(n2849));
  invx g2786(.A(n2851), .O(n2850));
  orx  g2787(.A(n3516), .B(n2852), .O(n2851));
  orx  g2788(.A(n2858), .B(n2853), .O(n2852));
  andx g2789(.A(n2854), .B(po12), .O(n2853));
  orx  g2790(.A(n2856), .B(n2855), .O(n2854));
  andx g2791(.A(n2976), .B(n2921), .O(n2855));
  andx g2792(.A(n2857), .B(n2975), .O(n2856));
  invx g2793(.A(n2921), .O(n2857));
  andx g2794(.A(n2980), .B(n158), .O(n2858));
  invx g2795(.A(n2860), .O(n2859));
  orx  g2796(.A(n2862), .B(n2861), .O(n2860));
  andx g2797(.A(n2864), .B(n3523), .O(n2861));
  invx g2798(.A(n2863), .O(n2862));
  orx  g2799(.A(n119), .B(n2864), .O(n2863));
  orx  g2800(.A(n2870), .B(n2865), .O(n2864));
  andx g2801(.A(n2866), .B(n2902), .O(n2865));
  orx  g2802(.A(n2868), .B(n2867), .O(n2866));
  andx g2803(.A(n2988), .B(n2919), .O(n2867));
  andx g2804(.A(n2869), .B(n2987), .O(n2868));
  invx g2805(.A(n2919), .O(n2869));
  andx g2806(.A(n2992), .B(n157), .O(n2870));
  invx g2807(.A(n2872), .O(n2871));
  orx  g2808(.A(n2874), .B(n2873), .O(n2872));
  andx g2809(.A(n2876), .B(n113), .O(n2873));
  invx g2810(.A(n2875), .O(n2874));
  orx  g2811(.A(n3524), .B(n2876), .O(n2875));
  orx  g2812(.A(n2882), .B(n2877), .O(n2876));
  andx g2813(.A(n2878), .B(po12), .O(n2877));
  orx  g2814(.A(n2880), .B(n2879), .O(n2878));
  andx g2815(.A(n3000), .B(n2917), .O(n2879));
  andx g2816(.A(n2881), .B(n2999), .O(n2880));
  invx g2817(.A(n2917), .O(n2881));
  andx g2818(.A(n3004), .B(n158), .O(n2882));
  invx g2819(.A(n2884), .O(n2883));
  orx  g2820(.A(n2886), .B(n2885), .O(n2884));
  andx g2821(.A(n2888), .B(n212), .O(n2885));
  invx g2822(.A(n2887), .O(n2886));
  orx  g2823(.A(n212), .B(n2888), .O(n2887));
  orx  g2824(.A(n2894), .B(n2889), .O(n2888));
  andx g2825(.A(n2890), .B(n2902), .O(n2889));
  orx  g2826(.A(n2892), .B(n2891), .O(n2890));
  andx g2827(.A(n3012), .B(n2915), .O(n2891));
  andx g2828(.A(n2893), .B(n3011), .O(n2892));
  invx g2829(.A(n2915), .O(n2893));
  andx g2830(.A(n3016), .B(n157), .O(n2894));
  invx g2831(.A(n2896), .O(n2895));
  andx g2832(.A(n2899), .B(n2897), .O(n2896));
  invx g2833(.A(n2898), .O(n2897));
  andx g2834(.A(n2900), .B(n211), .O(n2898));
  orx  g2835(.A(n208), .B(n2900), .O(n2899));
  orx  g2836(.A(n2904), .B(n2901), .O(n2900));
  andx g2837(.A(n2903), .B(po12), .O(n2901));
  invx g2838(.A(n157), .O(n2902));
  andx g2839(.A(n2909), .B(n2913), .O(n2903));
  andx g2840(.A(n3025), .B(n158), .O(n2904));
  orx  g2841(.A(n2907), .B(n2906), .O(n2905));
  invx g2842(.A(n3509), .O(n2906));
  andx g2843(.A(n3023), .B(n2908), .O(n2907));
  orx  g2844(.A(n2912), .B(n2909), .O(n2908));
  orx  g2845(.A(n2911), .B(n2910), .O(n2909));
  andx g2846(.A(n3025), .B(n215), .O(n2910));
  andx g2847(.A(pi19), .B(n3024), .O(n2911));
  invx g2848(.A(n2913), .O(n2912));
  orx  g2849(.A(n2914), .B(n3013), .O(n2913));
  andx g2850(.A(n3011), .B(n2915), .O(n2914));
  orx  g2851(.A(n2916), .B(n3001), .O(n2915));
  andx g2852(.A(n2999), .B(n2917), .O(n2916));
  orx  g2853(.A(n2918), .B(n2989), .O(n2917));
  andx g2854(.A(n2987), .B(n2919), .O(n2918));
  orx  g2855(.A(n2920), .B(n2977), .O(n2919));
  andx g2856(.A(n2975), .B(n2921), .O(n2920));
  orx  g2857(.A(n2922), .B(n2965), .O(n2921));
  andx g2858(.A(n2963), .B(n2923), .O(n2922));
  orx  g2859(.A(n2924), .B(n2953), .O(n2923));
  andx g2860(.A(n2951), .B(n2925), .O(n2924));
  orx  g2861(.A(n2926), .B(n2942), .O(n2925));
  andx g2862(.A(n2940), .B(n2927), .O(n2926));
  orx  g2863(.A(n2929), .B(n2928), .O(n2927));
  andx g2864(.A(n2936), .B(n218), .O(n2928));
  andx g2865(.A(n2931), .B(n65), .O(n2929));
  orx  g2866(.A(pi12), .B(n3500), .O(n2930));
  invx g2867(.A(n2932), .O(n2931));
  andx g2868(.A(n2934), .B(n2933), .O(n2932));
  orx  g2869(.A(n2936), .B(pi03), .O(n2933));
  invx g2870(.A(n2935), .O(n2934));
  andx g2871(.A(pi03), .B(n2936), .O(n2935));
  orx  g2872(.A(n2938), .B(n2937), .O(n2936));
  andx g2873(.A(n80), .B(n172), .O(n2937));
  andx g2874(.A(pi14), .B(n2939), .O(n2938));
  orx  g2875(.A(n3027), .B(n123), .O(n2939));
  invx g2876(.A(n2941), .O(n2940));
  orx  g2877(.A(n2943), .B(n2942), .O(n2941));
  andx g2878(.A(n2945), .B(n108), .O(n2942));
  invx g2879(.A(n2944), .O(n2943));
  orx  g2880(.A(n2945), .B(n137), .O(n2944));
  orx  g2881(.A(n2950), .B(n2946), .O(n2945));
  andx g2882(.A(n2947), .B(po14), .O(n2946));
  andx g2883(.A(n2949), .B(n2948), .O(n2947));
  orx  g2884(.A(n81), .B(n3050), .O(n2948));
  orx  g2885(.A(n80), .B(n3051), .O(n2949));
  andx g2886(.A(n3055), .B(n189), .O(n2950));
  invx g2887(.A(n2952), .O(n2951));
  orx  g2888(.A(n2954), .B(n2953), .O(n2952));
  andx g2889(.A(n2956), .B(n133), .O(n2953));
  invx g2890(.A(n2955), .O(n2954));
  orx  g2891(.A(n2956), .B(n135), .O(n2955));
  orx  g2892(.A(n2958), .B(n2957), .O(n2956));
  andx g2893(.A(n3064), .B(n189), .O(n2957));
  andx g2894(.A(n2959), .B(n172), .O(n2958));
  orx  g2895(.A(n2961), .B(n2960), .O(n2959));
  andx g2896(.A(n3060), .B(n3046), .O(n2960));
  andx g2897(.A(n2962), .B(n3059), .O(n2961));
  invx g2898(.A(n3046), .O(n2962));
  invx g2899(.A(n2964), .O(n2963));
  orx  g2900(.A(n2966), .B(n2965), .O(n2964));
  andx g2901(.A(n2968), .B(n131), .O(n2965));
  invx g2902(.A(n2967), .O(n2966));
  orx  g2903(.A(n2968), .B(n131), .O(n2967));
  orx  g2904(.A(n2970), .B(n2969), .O(n2968));
  andx g2905(.A(n3075), .B(n189), .O(n2969));
  andx g2906(.A(n2971), .B(po14), .O(n2970));
  orx  g2907(.A(n2973), .B(n2972), .O(n2971));
  andx g2908(.A(n3071), .B(n3044), .O(n2972));
  andx g2909(.A(n2974), .B(n3070), .O(n2973));
  invx g2910(.A(n3044), .O(n2974));
  invx g2911(.A(n2976), .O(n2975));
  orx  g2912(.A(n2978), .B(n2977), .O(n2976));
  andx g2913(.A(n2980), .B(n96), .O(n2977));
  invx g2914(.A(n2979), .O(n2978));
  orx  g2915(.A(n73), .B(n2980), .O(n2979));
  orx  g2916(.A(n2982), .B(n2981), .O(n2980));
  andx g2917(.A(n3087), .B(n189), .O(n2981));
  andx g2918(.A(n2983), .B(n172), .O(n2982));
  orx  g2919(.A(n2985), .B(n2984), .O(n2983));
  andx g2920(.A(n3083), .B(n3042), .O(n2984));
  andx g2921(.A(n2986), .B(n3082), .O(n2985));
  invx g2922(.A(n3042), .O(n2986));
  invx g2923(.A(n2988), .O(n2987));
  orx  g2924(.A(n2990), .B(n2989), .O(n2988));
  andx g2925(.A(n2992), .B(n3516), .O(n2989));
  invx g2926(.A(n2991), .O(n2990));
  orx  g2927(.A(n121), .B(n2992), .O(n2991));
  orx  g2928(.A(n2994), .B(n2993), .O(n2992));
  andx g2929(.A(n3099), .B(n189), .O(n2993));
  andx g2930(.A(n2995), .B(po14), .O(n2994));
  orx  g2931(.A(n2997), .B(n2996), .O(n2995));
  andx g2932(.A(n3095), .B(n3040), .O(n2996));
  andx g2933(.A(n2998), .B(n3094), .O(n2997));
  invx g2934(.A(n3040), .O(n2998));
  invx g2935(.A(n3000), .O(n2999));
  orx  g2936(.A(n3002), .B(n3001), .O(n3000));
  andx g2937(.A(n3004), .B(n116), .O(n3001));
  invx g2938(.A(n3003), .O(n3002));
  orx  g2939(.A(n119), .B(n3004), .O(n3003));
  orx  g2940(.A(n3006), .B(n3005), .O(n3004));
  andx g2941(.A(n3111), .B(n189), .O(n3005));
  andx g2942(.A(n3007), .B(n172), .O(n3006));
  orx  g2943(.A(n3009), .B(n3008), .O(n3007));
  andx g2944(.A(n3107), .B(n3038), .O(n3008));
  andx g2945(.A(n3010), .B(n3106), .O(n3009));
  invx g2946(.A(n3038), .O(n3010));
  invx g2947(.A(n3012), .O(n3011));
  orx  g2948(.A(n3014), .B(n3013), .O(n3012));
  andx g2949(.A(n3016), .B(n113), .O(n3013));
  invx g2950(.A(n3015), .O(n3014));
  orx  g2951(.A(n115), .B(n3016), .O(n3015));
  orx  g2952(.A(n3018), .B(n3017), .O(n3016));
  andx g2953(.A(n3123), .B(n3027), .O(n3017));
  andx g2954(.A(n3019), .B(po14), .O(n3018));
  orx  g2955(.A(n3021), .B(n3020), .O(n3019));
  andx g2956(.A(n3119), .B(n3036), .O(n3020));
  andx g2957(.A(n3022), .B(n3118), .O(n3021));
  invx g2958(.A(n3036), .O(n3022));
  orx  g2959(.A(pi19), .B(n3024), .O(n3023));
  invx g2960(.A(n3025), .O(n3024));
  orx  g2961(.A(n3028), .B(n3026), .O(n3025));
  andx g2962(.A(n3135), .B(n3027), .O(n3026));
  invx g2963(.A(po14), .O(n3027));
  andx g2964(.A(n3033), .B(n172), .O(n3028));
  orx  g2965(.A(n3031), .B(n3030), .O(n3029));
  andx g2966(.A(n3507), .B(n3135), .O(n3030));
  andx g2967(.A(n3032), .B(n3131), .O(n3031));
  andx g2968(.A(n3508), .B(n3034), .O(n3032));
  andx g2969(.A(n3130), .B(n3034), .O(n3033));
  orx  g2970(.A(n3035), .B(n3120), .O(n3034));
  andx g2971(.A(n3118), .B(n3036), .O(n3035));
  orx  g2972(.A(n3037), .B(n3108), .O(n3036));
  andx g2973(.A(n3106), .B(n3038), .O(n3037));
  orx  g2974(.A(n3039), .B(n3096), .O(n3038));
  andx g2975(.A(n3094), .B(n3040), .O(n3039));
  orx  g2976(.A(n3041), .B(n3084), .O(n3040));
  andx g2977(.A(n3082), .B(n3042), .O(n3041));
  orx  g2978(.A(n3043), .B(n3072), .O(n3042));
  andx g2979(.A(n3070), .B(n3044), .O(n3043));
  orx  g2980(.A(n3045), .B(n3061), .O(n3044));
  andx g2981(.A(n3059), .B(n3046), .O(n3045));
  orx  g2982(.A(n3048), .B(n3047), .O(n3046));
  andx g2983(.A(n3055), .B(n218), .O(n3047));
  andx g2984(.A(n3050), .B(n81), .O(n3048));
  orx  g2985(.A(pi14), .B(n123), .O(n3049));
  invx g2986(.A(n3051), .O(n3050));
  andx g2987(.A(n3053), .B(n3052), .O(n3051));
  orx  g2988(.A(n3055), .B(pi03), .O(n3052));
  invx g2989(.A(n3054), .O(n3053));
  andx g2990(.A(pi03), .B(n3055), .O(n3054));
  orx  g2991(.A(n3057), .B(n3056), .O(n3055));
  andx g2992(.A(n82), .B(n3139), .O(n3056));
  andx g2993(.A(pi16), .B(n3058), .O(n3057));
  orx  g2994(.A(n3137), .B(n91), .O(n3058));
  invx g2995(.A(n3060), .O(n3059));
  orx  g2996(.A(n3062), .B(n3061), .O(n3060));
  andx g2997(.A(n3064), .B(n137), .O(n3061));
  invx g2998(.A(n3063), .O(n3062));
  orx  g2999(.A(n3064), .B(n107), .O(n3063));
  orx  g3000(.A(n3069), .B(n3065), .O(n3064));
  andx g3001(.A(n3066), .B(n3139), .O(n3065));
  andx g3002(.A(n3068), .B(n3067), .O(n3066));
  orx  g3003(.A(n83), .B(n3158), .O(n3067));
  orx  g3004(.A(n82), .B(n3159), .O(n3068));
  andx g3005(.A(n3163), .B(n187), .O(n3069));
  invx g3006(.A(n3071), .O(n3070));
  orx  g3007(.A(n3073), .B(n3072), .O(n3071));
  andx g3008(.A(n3075), .B(n133), .O(n3072));
  invx g3009(.A(n3074), .O(n3073));
  orx  g3010(.A(n3075), .B(n104), .O(n3074));
  orx  g3011(.A(n3077), .B(n3076), .O(n3075));
  andx g3012(.A(n3172), .B(n187), .O(n3076));
  andx g3013(.A(n3078), .B(po16), .O(n3077));
  orx  g3014(.A(n3080), .B(n3079), .O(n3078));
  andx g3015(.A(n3168), .B(n3154), .O(n3079));
  andx g3016(.A(n3081), .B(n3167), .O(n3080));
  invx g3017(.A(n3154), .O(n3081));
  invx g3018(.A(n3083), .O(n3082));
  orx  g3019(.A(n3085), .B(n3084), .O(n3083));
  andx g3020(.A(n3087), .B(n3522), .O(n3084));
  invx g3021(.A(n3086), .O(n3085));
  orx  g3022(.A(n3087), .B(n131), .O(n3086));
  orx  g3023(.A(n3089), .B(n3088), .O(n3087));
  andx g3024(.A(n3183), .B(n187), .O(n3088));
  andx g3025(.A(n3090), .B(po16), .O(n3089));
  orx  g3026(.A(n3092), .B(n3091), .O(n3090));
  andx g3027(.A(n3179), .B(n3152), .O(n3091));
  andx g3028(.A(n3093), .B(n3178), .O(n3092));
  invx g3029(.A(n3152), .O(n3093));
  invx g3030(.A(n3095), .O(n3094));
  orx  g3031(.A(n3097), .B(n3096), .O(n3095));
  andx g3032(.A(n3099), .B(n129), .O(n3096));
  invx g3033(.A(n3098), .O(n3097));
  orx  g3034(.A(n95), .B(n3099), .O(n3098));
  orx  g3035(.A(n3101), .B(n3100), .O(n3099));
  andx g3036(.A(n3195), .B(n187), .O(n3100));
  andx g3037(.A(n3102), .B(po16), .O(n3101));
  orx  g3038(.A(n3104), .B(n3103), .O(n3102));
  andx g3039(.A(n3191), .B(n3150), .O(n3103));
  andx g3040(.A(n3105), .B(n3190), .O(n3104));
  invx g3041(.A(n3150), .O(n3105));
  invx g3042(.A(n3107), .O(n3106));
  orx  g3043(.A(n3109), .B(n3108), .O(n3107));
  andx g3044(.A(n3111), .B(n120), .O(n3108));
  invx g3045(.A(n3110), .O(n3109));
  orx  g3046(.A(n121), .B(n3111), .O(n3110));
  orx  g3047(.A(n3113), .B(n3112), .O(n3111));
  andx g3048(.A(n3207), .B(n187), .O(n3112));
  andx g3049(.A(n3114), .B(po16), .O(n3113));
  orx  g3050(.A(n3116), .B(n3115), .O(n3114));
  andx g3051(.A(n3203), .B(n3148), .O(n3115));
  andx g3052(.A(n3117), .B(n3202), .O(n3116));
  invx g3053(.A(n3148), .O(n3117));
  invx g3054(.A(n3119), .O(n3118));
  orx  g3055(.A(n3121), .B(n3120), .O(n3119));
  andx g3056(.A(n3123), .B(n119), .O(n3120));
  invx g3057(.A(n3122), .O(n3121));
  orx  g3058(.A(n119), .B(n3123), .O(n3122));
  orx  g3059(.A(n3125), .B(n3124), .O(n3123));
  andx g3060(.A(n3219), .B(n3137), .O(n3124));
  andx g3061(.A(n3126), .B(po16), .O(n3125));
  orx  g3062(.A(n3128), .B(n3127), .O(n3126));
  andx g3063(.A(n3215), .B(n3146), .O(n3127));
  andx g3064(.A(n3129), .B(n3214), .O(n3128));
  invx g3065(.A(n3146), .O(n3129));
  invx g3066(.A(n3131), .O(n3130));
  andx g3067(.A(n3134), .B(n3132), .O(n3131));
  invx g3068(.A(n3133), .O(n3132));
  andx g3069(.A(n3135), .B(n113), .O(n3133));
  orx  g3070(.A(n115), .B(n3135), .O(n3134));
  orx  g3071(.A(n3138), .B(n3136), .O(n3135));
  andx g3072(.A(n3231), .B(n3137), .O(n3136));
  invx g3073(.A(n3139), .O(n3137));
  andx g3074(.A(n3143), .B(po16), .O(n3138));
  orx  g3075(.A(n3141), .B(n3140), .O(n3139));
  andx g3076(.A(n3506), .B(n3231), .O(n3140));
  andx g3077(.A(n3142), .B(n3227), .O(n3141));
  andx g3078(.A(n3507), .B(n3144), .O(n3142));
  andx g3079(.A(n3226), .B(n3144), .O(n3143));
  orx  g3080(.A(n3145), .B(n3216), .O(n3144));
  andx g3081(.A(n3214), .B(n3146), .O(n3145));
  orx  g3082(.A(n3147), .B(n3204), .O(n3146));
  andx g3083(.A(n3202), .B(n3148), .O(n3147));
  orx  g3084(.A(n3149), .B(n3192), .O(n3148));
  andx g3085(.A(n3190), .B(n3150), .O(n3149));
  orx  g3086(.A(n3151), .B(n3180), .O(n3150));
  andx g3087(.A(n3178), .B(n3152), .O(n3151));
  orx  g3088(.A(n3153), .B(n3169), .O(n3152));
  andx g3089(.A(n3167), .B(n3154), .O(n3153));
  orx  g3090(.A(n3156), .B(n3155), .O(n3154));
  andx g3091(.A(n3163), .B(n219), .O(n3155));
  andx g3092(.A(n3158), .B(n83), .O(n3156));
  orx  g3093(.A(pi16), .B(n124), .O(n3157));
  invx g3094(.A(n3159), .O(n3158));
  andx g3095(.A(n3161), .B(n3160), .O(n3159));
  orx  g3096(.A(n3163), .B(pi03), .O(n3160));
  invx g3097(.A(n3162), .O(n3161));
  andx g3098(.A(pi03), .B(n3163), .O(n3162));
  orx  g3099(.A(n3165), .B(n3164), .O(n3163));
  andx g3100(.A(po18), .B(n84), .O(n3164));
  andx g3101(.A(pi18), .B(n3166), .O(n3165));
  orx  g3102(.A(n123), .B(n166), .O(n3166));
  invx g3103(.A(n3168), .O(n3167));
  orx  g3104(.A(n3170), .B(n3169), .O(n3168));
  andx g3105(.A(n3172), .B(n139), .O(n3169));
  invx g3106(.A(n3171), .O(n3170));
  orx  g3107(.A(n3172), .B(n137), .O(n3171));
  orx  g3108(.A(n3177), .B(n3173), .O(n3172));
  andx g3109(.A(n3174), .B(po18), .O(n3173));
  andx g3110(.A(n3176), .B(n3175), .O(n3174));
  orx  g3111(.A(n85), .B(n3256), .O(n3175));
  orx  g3112(.A(n84), .B(n3257), .O(n3176));
  andx g3113(.A(n3261), .B(n166), .O(n3177));
  invx g3114(.A(n3179), .O(n3178));
  orx  g3115(.A(n3181), .B(n3180), .O(n3179));
  andx g3116(.A(n3183), .B(n135), .O(n3180));
  invx g3117(.A(n3182), .O(n3181));
  orx  g3118(.A(n3183), .B(n133), .O(n3182));
  orx  g3119(.A(n3189), .B(n3184), .O(n3183));
  andx g3120(.A(n3185), .B(po18), .O(n3184));
  orx  g3121(.A(n3187), .B(n3186), .O(n3185));
  andx g3122(.A(n3266), .B(n3252), .O(n3186));
  andx g3123(.A(n3188), .B(n3265), .O(n3187));
  invx g3124(.A(n3252), .O(n3188));
  andx g3125(.A(n3270), .B(n166), .O(n3189));
  invx g3126(.A(n3191), .O(n3190));
  orx  g3127(.A(n3193), .B(n3192), .O(n3191));
  andx g3128(.A(n3195), .B(n132), .O(n3192));
  invx g3129(.A(n3194), .O(n3193));
  orx  g3130(.A(n3195), .B(n131), .O(n3194));
  orx  g3131(.A(n3201), .B(n3196), .O(n3195));
  andx g3132(.A(n3197), .B(po18), .O(n3196));
  orx  g3133(.A(n3199), .B(n3198), .O(n3197));
  andx g3134(.A(n3277), .B(n3250), .O(n3198));
  andx g3135(.A(n3200), .B(n3276), .O(n3199));
  invx g3136(.A(n3250), .O(n3200));
  andx g3137(.A(n3281), .B(n166), .O(n3201));
  invx g3138(.A(n3203), .O(n3202));
  orx  g3139(.A(n3205), .B(n3204), .O(n3203));
  andx g3140(.A(n3207), .B(n73), .O(n3204));
  invx g3141(.A(n3206), .O(n3205));
  orx  g3142(.A(n127), .B(n3207), .O(n3206));
  orx  g3143(.A(n3213), .B(n3208), .O(n3207));
  andx g3144(.A(n3209), .B(po18), .O(n3208));
  orx  g3145(.A(n3211), .B(n3210), .O(n3209));
  andx g3146(.A(n3289), .B(n3248), .O(n3210));
  andx g3147(.A(n3212), .B(n3288), .O(n3211));
  invx g3148(.A(n3248), .O(n3212));
  andx g3149(.A(n3293), .B(n166), .O(n3213));
  invx g3150(.A(n3215), .O(n3214));
  orx  g3151(.A(n3217), .B(n3216), .O(n3215));
  andx g3152(.A(n3219), .B(n94), .O(n3216));
  invx g3153(.A(n3218), .O(n3217));
  orx  g3154(.A(n121), .B(n3219), .O(n3218));
  orx  g3155(.A(n3225), .B(n3220), .O(n3219));
  andx g3156(.A(n3221), .B(po18), .O(n3220));
  orx  g3157(.A(n3223), .B(n3222), .O(n3221));
  andx g3158(.A(n3300), .B(n3246), .O(n3222));
  andx g3159(.A(n3224), .B(n3299), .O(n3223));
  invx g3160(.A(n3246), .O(n3224));
  andx g3161(.A(n3304), .B(n3236), .O(n3225));
  invx g3162(.A(n3227), .O(n3226));
  andx g3163(.A(n3230), .B(n3228), .O(n3227));
  invx g3164(.A(n3229), .O(n3228));
  andx g3165(.A(n3231), .B(n117), .O(n3229));
  orx  g3166(.A(n90), .B(n3231), .O(n3230));
  orx  g3167(.A(n3235), .B(n3232), .O(n3231));
  andx g3168(.A(n3234), .B(po18), .O(n3232));
  invx g3169(.A(n3236), .O(po18));
  andx g3170(.A(n3240), .B(n3244), .O(n3234));
  andx g3171(.A(n3313), .B(n3236), .O(n3235));
  orx  g3172(.A(n3238), .B(n3237), .O(n3236));
  invx g3173(.A(n3506), .O(n3237));
  andx g3174(.A(n3311), .B(n3239), .O(n3238));
  orx  g3175(.A(n3243), .B(n3240), .O(n3239));
  orx  g3176(.A(n3242), .B(n3241), .O(n3240));
  andx g3177(.A(n3313), .B(n120), .O(n3241));
  andx g3178(.A(pi13), .B(n3312), .O(n3242));
  invx g3179(.A(n3244), .O(n3243));
  orx  g3180(.A(n3245), .B(n3301), .O(n3244));
  andx g3181(.A(n3299), .B(n3246), .O(n3245));
  orx  g3182(.A(n3247), .B(n3290), .O(n3246));
  andx g3183(.A(n3288), .B(n3248), .O(n3247));
  orx  g3184(.A(n3249), .B(n3278), .O(n3248));
  andx g3185(.A(n3276), .B(n3250), .O(n3249));
  orx  g3186(.A(n3251), .B(n3267), .O(n3250));
  andx g3187(.A(n3265), .B(n3252), .O(n3251));
  orx  g3188(.A(n3254), .B(n3253), .O(n3252));
  andx g3189(.A(n3261), .B(n164), .O(n3253));
  andx g3190(.A(n3256), .B(n85), .O(n3254));
  orx  g3191(.A(pi18), .B(n124), .O(n3255));
  invx g3192(.A(n3257), .O(n3256));
  andx g3193(.A(n3259), .B(n3258), .O(n3257));
  orx  g3194(.A(n3261), .B(pi03), .O(n3258));
  invx g3195(.A(n3260), .O(n3259));
  andx g3196(.A(pi03), .B(n3261), .O(n3260));
  orx  g3197(.A(n3263), .B(n3262), .O(n3261));
  andx g3198(.A(n86), .B(po20), .O(n3262));
  andx g3199(.A(pi20), .B(n3264), .O(n3263));
  orx  g3200(.A(n3315), .B(n91), .O(n3264));
  invx g3201(.A(n3266), .O(n3265));
  orx  g3202(.A(n3268), .B(n3267), .O(n3266));
  andx g3203(.A(n3270), .B(n137), .O(n3267));
  invx g3204(.A(n3269), .O(n3268));
  orx  g3205(.A(n3270), .B(n105), .O(n3269));
  orx  g3206(.A(n3275), .B(n3271), .O(n3270));
  andx g3207(.A(n3272), .B(po20), .O(n3271));
  andx g3208(.A(n3274), .B(n3273), .O(n3272));
  orx  g3209(.A(n87), .B(n3349), .O(n3273));
  orx  g3210(.A(n86), .B(n3350), .O(n3274));
  andx g3211(.A(n3354), .B(n3315), .O(n3275));
  invx g3212(.A(n3277), .O(n3276));
  orx  g3213(.A(n3279), .B(n3278), .O(n3277));
  andx g3214(.A(n3281), .B(n3517), .O(n3278));
  invx g3215(.A(n3280), .O(n3279));
  orx  g3216(.A(n3281), .B(n103), .O(n3280));
  orx  g3217(.A(n3283), .B(n3282), .O(n3281));
  andx g3218(.A(n3363), .B(n3315), .O(n3282));
  andx g3219(.A(n3284), .B(po20), .O(n3283));
  orx  g3220(.A(n3286), .B(n3285), .O(n3284));
  andx g3221(.A(n3359), .B(n3345), .O(n3285));
  andx g3222(.A(n3287), .B(n3358), .O(n3286));
  invx g3223(.A(n3345), .O(n3287));
  invx g3224(.A(n3289), .O(n3288));
  orx  g3225(.A(n3291), .B(n3290), .O(n3289));
  andx g3226(.A(n3293), .B(n132), .O(n3290));
  invx g3227(.A(n3292), .O(n3291));
  orx  g3228(.A(n3293), .B(n3522), .O(n3292));
  orx  g3229(.A(n3298), .B(n3294), .O(n3293));
  andx g3230(.A(n3295), .B(po20), .O(n3294));
  andx g3231(.A(n3297), .B(n3296), .O(n3295));
  orx  g3232(.A(n3328), .B(n3343), .O(n3296));
  invx g3233(.A(n3327), .O(n3297));
  andx g3234(.A(n3332), .B(n3315), .O(n3298));
  invx g3235(.A(n3300), .O(n3299));
  orx  g3236(.A(n3302), .B(n3301), .O(n3300));
  andx g3237(.A(n3304), .B(n129), .O(n3301));
  invx g3238(.A(n3303), .O(n3302));
  orx  g3239(.A(n127), .B(n3304), .O(n3303));
  orx  g3240(.A(n3306), .B(n3305), .O(n3304));
  andx g3241(.A(n3378), .B(n3315), .O(n3305));
  andx g3242(.A(n3307), .B(po20), .O(n3306));
  orx  g3243(.A(n3309), .B(n3308), .O(n3307));
  andx g3244(.A(n3374), .B(n3325), .O(n3308));
  andx g3245(.A(n3310), .B(n3373), .O(n3309));
  invx g3246(.A(n3325), .O(n3310));
  orx  g3247(.A(pi13), .B(n3312), .O(n3311));
  invx g3248(.A(n3313), .O(n3312));
  orx  g3249(.A(n3316), .B(n3314), .O(n3313));
  andx g3250(.A(n3391), .B(n3315), .O(n3314));
  invx g3251(.A(po20), .O(n3315));
  andx g3252(.A(n3322), .B(po20), .O(n3316));
  orx  g3253(.A(n3319), .B(n3318), .O(n3317));
  andx g3254(.A(n3504), .B(n3391), .O(n3318));
  andx g3255(.A(n3321), .B(n3320), .O(n3319));
  invx g3256(.A(n3387), .O(n3320));
  andx g3257(.A(n3505), .B(n3323), .O(n3321));
  andx g3258(.A(n3387), .B(n3323), .O(n3322));
  orx  g3259(.A(n3324), .B(n3375), .O(n3323));
  andx g3260(.A(n3373), .B(n3325), .O(n3324));
  orx  g3261(.A(n3327), .B(n3326), .O(n3325));
  andx g3262(.A(n3332), .B(n135), .O(n3326));
  andx g3263(.A(n3343), .B(n3328), .O(n3327));
  orx  g3264(.A(n3331), .B(n3329), .O(n3328));
  invx g3265(.A(n3330), .O(n3329));
  orx  g3266(.A(n3332), .B(pi07), .O(n3330));
  andx g3267(.A(pi07), .B(n3332), .O(n3331));
  orx  g3268(.A(n3336), .B(n3333), .O(n3332));
  andx g3269(.A(n3427), .B(n3334), .O(n3333));
  orx  g3270(.A(n3393), .B(n3335), .O(n3334));
  andx g3271(.A(n3339), .B(n107), .O(n3335));
  andx g3272(.A(n3337), .B(po22), .O(n3336));
  andx g3273(.A(n3339), .B(n3338), .O(n3337));
  invx g3274(.A(n3413), .O(n3338));
  orx  g3275(.A(n3340), .B(n3414), .O(n3339));
  andx g3276(.A(n3341), .B(n3425), .O(n3340));
  orx  g3277(.A(pi05), .B(n3342), .O(n3341));
  invx g3278(.A(n3427), .O(n3342));
  orx  g3279(.A(n3344), .B(n3360), .O(n3343));
  andx g3280(.A(n3358), .B(n3345), .O(n3344));
  orx  g3281(.A(n3347), .B(n3346), .O(n3345));
  andx g3282(.A(n3354), .B(n216), .O(n3346));
  andx g3283(.A(n3349), .B(n87), .O(n3347));
  orx  g3284(.A(pi20), .B(n126), .O(n3348));
  invx g3285(.A(n3350), .O(n3349));
  andx g3286(.A(n3352), .B(n3351), .O(n3350));
  orx  g3287(.A(n3354), .B(pi03), .O(n3351));
  invx g3288(.A(n3353), .O(n3352));
  andx g3289(.A(pi03), .B(n3354), .O(n3353));
  orx  g3290(.A(n3356), .B(n3355), .O(n3354));
  andx g3291(.A(po22), .B(n3419), .O(n3355));
  andx g3292(.A(pi22), .B(n3357), .O(n3356));
  orx  g3293(.A(n124), .B(n3393), .O(n3357));
  invx g3294(.A(n3359), .O(n3358));
  orx  g3295(.A(n3361), .B(n3360), .O(n3359));
  andx g3296(.A(n3363), .B(n3518), .O(n3360));
  invx g3297(.A(n3362), .O(n3361));
  orx  g3298(.A(n3363), .B(n3518), .O(n3362));
  orx  g3299(.A(n3370), .B(n3364), .O(n3363));
  andx g3300(.A(n3366), .B(n3365), .O(n3364));
  invx g3301(.A(n3421), .O(n3365));
  andx g3302(.A(po22), .B(n3367), .O(n3366));
  orx  g3303(.A(n3369), .B(n3368), .O(n3367));
  andx g3304(.A(n3419), .B(n217), .O(n3368));
  andx g3305(.A(pi03), .B(n3420), .O(n3369));
  andx g3306(.A(n3371), .B(n3421), .O(n3370));
  orx  g3307(.A(n3372), .B(n3393), .O(n3371));
  orx  g3308(.A(n3415), .B(n3418), .O(n3372));
  invx g3309(.A(n3374), .O(n3373));
  orx  g3310(.A(n3376), .B(n3375), .O(n3374));
  andx g3311(.A(n3378), .B(n132), .O(n3375));
  invx g3312(.A(n3377), .O(n3376));
  orx  g3313(.A(n3378), .B(n132), .O(n3377));
  orx  g3314(.A(n3386), .B(n3379), .O(n3378));
  andx g3315(.A(n3380), .B(po22), .O(n3379));
  andx g3316(.A(n3383), .B(n3381), .O(n3380));
  invx g3317(.A(n3382), .O(n3381));
  andx g3318(.A(n3412), .B(n3384), .O(n3382));
  orx  g3319(.A(n3384), .B(n3412), .O(n3383));
  andx g3320(.A(n3402), .B(n3385), .O(n3384));
  invx g3321(.A(n3400), .O(n3385));
  andx g3322(.A(n3403), .B(n3393), .O(n3386));
  andx g3323(.A(n3389), .B(n3388), .O(n3387));
  orx  g3324(.A(n3391), .B(pi11), .O(n3388));
  invx g3325(.A(n3390), .O(n3389));
  andx g3326(.A(pi11), .B(n3391), .O(n3390));
  orx  g3327(.A(n3398), .B(n3392), .O(n3391));
  andx g3328(.A(n3438), .B(n3393), .O(n3392));
  invx g3329(.A(po22), .O(n3393));
  andx g3330(.A(n3395), .B(n3504), .O(po22));
  orx  g3331(.A(n3437), .B(n3396), .O(n3395));
  andx g3332(.A(n3399), .B(n3397), .O(n3396));
  orx  g3333(.A(n3438), .B(n132), .O(n3397));
  andx g3334(.A(n3437), .B(n3399), .O(n3398));
  orx  g3335(.A(n3401), .B(n3400), .O(n3399));
  andx g3336(.A(n133), .B(n3403), .O(n3400));
  andx g3337(.A(n3412), .B(n3402), .O(n3401));
  orx  g3338(.A(n104), .B(n3403), .O(n3402));
  orx  g3339(.A(n3407), .B(n3404), .O(n3403));
  andx g3340(.A(n3463), .B(n3405), .O(n3404));
  orx  g3341(.A(n3440), .B(n3406), .O(n3405));
  andx g3342(.A(n3408), .B(n71), .O(n3406));
  andx g3343(.A(n3410), .B(n3408), .O(n3407));
  orx  g3344(.A(n3409), .B(n3450), .O(n3408));
  andx g3345(.A(pi05), .B(n3449), .O(n3409));
  invx g3346(.A(n3411), .O(n3410));
  orx  g3347(.A(n3440), .B(n3448), .O(n3411));
  orx  g3348(.A(n3413), .B(n3426), .O(n3412));
  andx g3349(.A(n3425), .B(n3414), .O(n3413));
  orx  g3350(.A(n3416), .B(n3415), .O(n3414));
  andx g3351(.A(n218), .B(n3420), .O(n3415));
  andx g3352(.A(n3421), .B(n3417), .O(n3416));
  invx g3353(.A(n3418), .O(n3417));
  andx g3354(.A(pi03), .B(n3419), .O(n3418));
  invx g3355(.A(n3420), .O(n3419));
  orx  g3356(.A(pi22), .B(n126), .O(n3420));
  orx  g3357(.A(n3423), .B(n3422), .O(n3421));
  andx g3358(.A(n3455), .B(po24), .O(n3422));
  andx g3359(.A(pi24), .B(n3424), .O(n3423));
  orx  g3360(.A(n3440), .B(n91), .O(n3424));
  orx  g3361(.A(n138), .B(n3427), .O(n3425));
  andx g3362(.A(n3427), .B(n3518), .O(n3426));
  orx  g3363(.A(n3434), .B(n3428), .O(n3427));
  andx g3364(.A(n3430), .B(n3429), .O(n3428));
  invx g3365(.A(n3457), .O(n3429));
  andx g3366(.A(n3431), .B(po24), .O(n3430));
  orx  g3367(.A(n3433), .B(n3432), .O(n3431));
  andx g3368(.A(n3455), .B(n217), .O(n3432));
  andx g3369(.A(pi03), .B(n3456), .O(n3433));
  andx g3370(.A(n3435), .B(n3457), .O(n3434));
  orx  g3371(.A(n3440), .B(n3436), .O(n3435));
  orx  g3372(.A(n3451), .B(n3454), .O(n3436));
  andx g3373(.A(n130), .B(n3438), .O(n3437));
  orx  g3374(.A(n3446), .B(n3439), .O(n3438));
  andx g3375(.A(n3470), .B(n3440), .O(n3439));
  invx g3376(.A(po24), .O(n3440));
  orx  g3377(.A(n3443), .B(n3442), .O(po24));
  andx g3378(.A(n3502), .B(n3470), .O(n3442));
  andx g3379(.A(n3444), .B(n3503), .O(n3443));
  andx g3380(.A(n3447), .B(n3445), .O(n3444));
  orx  g3381(.A(n3470), .B(n103), .O(n3445));
  andx g3382(.A(n3469), .B(n3447), .O(n3446));
  orx  g3383(.A(n3448), .B(n3462), .O(n3447));
  andx g3384(.A(n3450), .B(n3449), .O(n3448));
  orx  g3385(.A(n107), .B(n3463), .O(n3449));
  orx  g3386(.A(n3452), .B(n3451), .O(n3450));
  andx g3387(.A(n217), .B(n3456), .O(n3451));
  andx g3388(.A(n3457), .B(n3453), .O(n3452));
  invx g3389(.A(n3454), .O(n3453));
  andx g3390(.A(pi03), .B(n3455), .O(n3454));
  invx g3391(.A(n3456), .O(n3455));
  orx  g3392(.A(pi24), .B(n125), .O(n3456));
  orx  g3393(.A(n3460), .B(n3458), .O(n3457));
  andx g3394(.A(n3459), .B(po26), .O(n3458));
  invx g3395(.A(n3483), .O(n3459));
  andx g3396(.A(pi26), .B(n3461), .O(n3460));
  orx  g3397(.A(n3473), .B(n125), .O(n3461));
  andx g3398(.A(n3463), .B(n108), .O(n3462));
  orx  g3399(.A(n3467), .B(n3464), .O(n3463));
  andx g3400(.A(n3465), .B(n3485), .O(n3464));
  andx g3401(.A(n3466), .B(po26), .O(n3465));
  andx g3402(.A(n3483), .B(pi03), .O(n3466));
  andx g3403(.A(n3468), .B(n3484), .O(n3467));
  orx  g3404(.A(n3480), .B(n3473), .O(n3468));
  andx g3405(.A(n3470), .B(n135), .O(n3469));
  andx g3406(.A(n3471), .B(n3487), .O(n3470));
  orx  g3407(.A(n3473), .B(n3472), .O(n3471));
  andx g3408(.A(n71), .B(n3479), .O(n3472));
  invx g3409(.A(po26), .O(n3473));
  orx  g3410(.A(n3476), .B(n3475), .O(po26));
  andx g3411(.A(n93), .B(n3479), .O(n3475));
  andx g3412(.A(n3487), .B(n3477), .O(n3476));
  orx  g3413(.A(n3478), .B(n93), .O(n3477));
  andx g3414(.A(n3502), .B(n3479), .O(n3478));
  orx  g3415(.A(n3481), .B(n3480), .O(n3479));
  andx g3416(.A(n216), .B(n3483), .O(n3480));
  andx g3417(.A(n3484), .B(n3482), .O(n3481));
  orx  g3418(.A(n3483), .B(n164), .O(n3482));
  orx  g3419(.A(pi26), .B(n123), .O(n3483));
  invx g3420(.A(n3485), .O(n3484));
  orx  g3421(.A(n3486), .B(n3521), .O(n3485));
  andx g3422(.A(po28), .B(pi01), .O(n3486));
  invx g3423(.A(n3488), .O(n3487));
  orx  g3424(.A(n3489), .B(n3494), .O(n3488));
  andx g3425(.A(po28), .B(n3519), .O(n3489));
  andx g3426(.A(n3491), .B(n93), .O(po28));
  invx g3427(.A(n3492), .O(n3491));
  andx g3428(.A(n3519), .B(n3493), .O(n3492));
  orx  g3429(.A(n3520), .B(n3494), .O(n3493));
  orx  g3430(.A(n3496), .B(n3495), .O(n3494));
  invx g3431(.A(pi30), .O(n3495));
  andx g3432(.A(po30), .B(pi01), .O(n3496));
  andx g3433(.A(n93), .B(n3498), .O(po30));
  andx g3434(.A(n219), .B(n3499), .O(n3498));
  orx  g3435(.A(n126), .B(pi30), .O(n3499));
  invx g3436(.A(pi01), .O(n3500));
  andx g3437(.A(n138), .B(n3502), .O(n3501));
  andx g3438(.A(n135), .B(n3503), .O(n3502));
  andx g3439(.A(n132), .B(n3504), .O(n3503));
  andx g3440(.A(n127), .B(n3505), .O(n3504));
  andx g3441(.A(n72), .B(n3506), .O(n3505));
  andx g3442(.A(n116), .B(n3507), .O(n3506));
  andx g3443(.A(n113), .B(n3508), .O(n3507));
  andx g3444(.A(n213), .B(n3509), .O(n3508));
  andx g3445(.A(n211), .B(n3510), .O(n3509));
  andx g3446(.A(n198), .B(n3511), .O(n3510));
  andx g3447(.A(n143), .B(n3512), .O(n3511));
  andx g3448(.A(n141), .B(n3513), .O(n3512));
  andx g3449(.A(n3514), .B(n3529), .O(n3513));
  invx g3450(.A(pi31), .O(n3514));
  invx g3451(.A(pi19), .O(n3515));
  invx g3452(.A(pi13), .O(n3516));
  invx g3453(.A(pi07), .O(n3517));
  invx g3454(.A(pi05), .O(n3518));
  orx  g3455(.A(pi03), .B(n3520), .O(n3519));
  andx g3456(.A(n3521), .B(pi01), .O(n3520));
  invx g3457(.A(pi28), .O(n3521));
  invx g3458(.A(pi09), .O(n3522));
  invx g3459(.A(pi15), .O(n3523));
  invx g3460(.A(pi17), .O(n3524));
  invx g3461(.A(pi21), .O(n3525));
  invx g3462(.A(pi23), .O(n3526));
  invx g3463(.A(pi25), .O(n3527));
  invx g3464(.A(pi27), .O(n3528));
  invx g3465(.A(pi29), .O(n3529));
endmodule


