// Benchmark "REVX" written by ABC on Wed Oct 16 00:55:51 2013

module REVX ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24;
  wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n131, n132, n133, n135, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
    n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
    n682, n683, n684, n685, n686, n687, n691, n692, n693, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n947, n948, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1267, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
    n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2155, n2156, n2157, n2158, n2161, n2162, n2164, n2167,
    n2168, n2169, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2392, n2393, n2394,
    n2395, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2432, n2439, n2450, n2452, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2523, n2524, n2525, n2526, n2527, n2530, n2531, n2532, n2535,
    n2536, n2537, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
    n2684, n2687, n2688, n2694, n2695, n2696, n2697, n2702, n2703, n2704,
    n2705, n2722, n2723, n2724, n2730, n2732, n2734, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2756, n2757,
    n2758, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816, n2818, n2821, n2827, n2828,
    n2829, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2879, n2880,
    n2883, n2884, n2888, n2889, n2890, n2891, n2895, n2896, n2899, n2900,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2989, n2990, n2994, n2996, n3001, n3005, n3006, n3007, n3008,
    n3011, n3013, n3014, n3015, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3027, n3028, n3031, n3033, n3034, n3035, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3091,
    n3092, n3096, n3097, n3098, n3099, n3100, n3103, n3104, n3105, n3107,
    n3108, n3113, n3114, n3119, n3120, n3121, n3122, n3126, n3127, n3128,
    n3129, n3131, n3132, n3136, n3137, n3138, n3139, n3144, n3145, n3151,
    n3152, n3153, n3154, n3156, n3157, n3158, n3159, n3160, n3161, n3166,
    n3167, n3168, n3169, n3170, n3171, n3175, n3179, n3180, n3181, n3182,
    n3183, n3185, n3194, n3200, n3201, n3202, n3205, n3206, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3292,
    n3293, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3345, n3346, n3347, n3348, n3349, n3353,
    n3354, n3355, n3357, n3358, n3359, n3360, n3361, n3363, n3366, n3367,
    n3368, n3369, n3370, n3372, n3373, n3374, n3379, n3380, n3383, n3384,
    n3388, n3389, n3390, n3391, n3395, n3396, n3397, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
    n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
    n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
    n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3566, n3567, n3568, n3569, n3570, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3582, n3585, n3586, n3587,
    n3588, n3589, n3590, n3591, n3593, n3596, n3597, n3603, n3604, n3605,
    n3606, n3607, n3608, n3612, n3614, n3615, n3616, n3619, n3620, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
    n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
    n3662, n3663, n3664, n3668, n3670, n3671, n3674, n3675, n3676, n3678,
    n3681, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
    n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
    n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
    n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
    n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4039,
    n4043, n4044, n4047, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4100, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4466, n4468, n4469, n4470, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4709, n4710,
    n4716, n4717, n4718, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
    n4727, n4728, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
    n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4980, n4983,
    n4984, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
    n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5085, n5086, n5087,
    n5088, n5098, n5099, n5100, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5131, n5132, n5133, n5134, n5138, n5139, n5143, n5144,
    n5145, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5381,
    n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398, n5400, n5401, n5402, n5403,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5460, n5461, n5462, n5466, n5467,
    n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
    n5478, n5488, n5489, n5490, n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
    n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
    n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
    n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5830,
    n5831, n5832, n5833, n5834, n5835, n5838, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5851, n5852, n5853, n5855, n5856, n5858, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5878, n5888, n5889, n5890, n5894, n5895,
    n5896, n5897, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6045, n6046, n6047, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
    n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6129, n6130, n6131, n6132, n6133, n6143, n6144, n6145, n6146,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6231,
    n6232, n6233, n6234, n6236, n6237, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6273,
    n6274, n6275, n6279, n6280, n6281, n6282, n6292, n6293, n6294, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6320, n6321, n6322, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
    n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
    n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
    n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6572, n6573,
    n6576, n6577, n6578, n6579, n6580, n6582, n6583, n6584, n6585, n6586,
    n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6619, n6620, n6621, n6622, n6626, n6627, n6628,
    n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
    n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
    n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
    n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
    n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
    n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6855, n6856,
    n6857, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
    n6888, n6889, n6890, n6891, n6894, n6895, n6896, n6897, n6898, n6899,
    n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
    n6911, n6912, n6913, n6914, n6916, n6917, n6918, n6920, n6921, n6924,
    n6925, n6926, n6927, n6929, n6930, n6931, n6932, n6933, n6936, n6937,
    n6940, n6941, n6942, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
    n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7030, n7031, n7032, n7033, n7034,
    n7035, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
    n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
    n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7257, n7259, n7261,
    n7262, n7263, n7264, n7266, n7267, n7268, n7269, n7270, n7273, n7276,
    n7277, n7278, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
    n7300, n7304, n7305, n7306, n7308, n7310, n7312, n7314, n7315, n7323,
    n7324, n7325, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7381,
    n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7397, n7398,
    n7399, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
    n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
    n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
    n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
    n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7624, n7625, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7644, n7646, n7652, n7653, n7654, n7655,
    n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
    n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
    n7697, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7712, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
    n7736, n7737, n7738, n7740, n7742, n7743, n7744, n7745, n7746, n7747,
    n7756, n7757, n7758, n7759, n7760, n7761, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7821, n7822, n7823, n7825,
    n7826, n7827, n7828, n7829, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8315, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
    n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
    n8350, n8351, n8352, n8353, n8361, n8362, n8363, n8364, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
    n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
    n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
    n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
    n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8506, n8507, n8508, n8510, n8511, n8512, n8513, n8514, n8515,
    n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
    n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
    n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
    n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
    n8656, n8657, n8658, n8663, n8664, n8665, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8836, n8837, n8838,
    n8839, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
    n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
    n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
    n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
    n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
    n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
    n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
    n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
    n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9060, n9061, n9062, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
    n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
    n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
    n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
    n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
    n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
    n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
    n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
    n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
    n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
    n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
    n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
    n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9710, n9711, n9712,
    n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
    n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
    n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
    n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
    n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
    n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
    n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
    n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
    n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
    n10024, n10033, n10034, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10072,
    n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10152, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10293, n10294, n10295, n10296,
    n10297, n10298, n10300, n10302, n10303, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
    n10320, n10321, n10322, n10323, n10324, n10329, n10330, n10332, n10333,
    n10334, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
    n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
    n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10370, n10371,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
    n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
    n10488, n10489, n10490, n10491, n10495, n10496, n10497, n10498, n10499,
    n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
    n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10703, n10704, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
    n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
    n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10844, n10848,
    n10849, n10850, n10851, n10852, n10854, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
    n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
    n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
    n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
    n11100, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
    n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
    n11147, n11150, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11164, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
    n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
    n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
    n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
    n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
    n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
    n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
    n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
    n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
    n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
    n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
    n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
    n11418, n11419, n11420, n11421, n11423, n11424, n11425, n11426, n11427,
    n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
    n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
    n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
    n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11463, n11464,
    n11465, n11466, n11467, n11471, n11474, n11475, n11477, n11480, n11481,
    n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11496, n11497, n11498, n11499, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
    n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
    n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
    n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
    n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
    n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
    n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
    n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
    n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759, n11761, n11762, n11763,
    n11764, n11765, n11766, n11767, n11768, n11769, n11772, n11775, n11776,
    n11777, n11778, n11779, n11780, n11781, n11782, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
    n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
    n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
    n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
    n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
    n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
    n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
    n12036, n12037, n12038, n12039, n12040, n12042, n12043, n12044, n12045,
    n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12056,
    n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
    n12069, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
    n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
    n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
    n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
    n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
    n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
    n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
    n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
    n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
    n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
    n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
    n12338, n12341, n12342, n12344, n12348, n12350, n12351, n12352, n12353,
    n12354, n12355, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
    n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
    n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
    n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
    n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
    n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
    n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
    n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
    n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12559, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12572, n12578, n12579, n12580, n12581, n12582,
    n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
    n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
    n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
    n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
    n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
    n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
    n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
    n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
    n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
    n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
    n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
    n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
    n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
    n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
    n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
    n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
    n12745, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
    n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
    n12764, n12765, n12766, n12767, n12768, n12769, n12782, n12783, n12786,
    n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
    n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
    n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
    n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
    n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
    n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
    n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
    n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
    n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
    n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
    n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
    n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
    n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
    n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
    n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
    n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
    n12940, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
    n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
    n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
    n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
    n12977, n12978, n12979, n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12999, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
    n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
    n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
    n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
    n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
    n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
    n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
    n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
    n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
    n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
    n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13145,
    n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
    n13164, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13189, n13190, n13191, n13192, n13193,
    n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
    n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
    n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
    n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
    n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
    n13312, n13313, n13314, n13315, n13316, n13317, n13320, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
    n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
    n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
    n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13436, n13437, n13438, n13439, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13471, n13474,
    n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
    n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
    n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
    n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
    n13556, n13557, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
    n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13585,
    n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
    n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
    n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
    n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
    n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13679, n13680, n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13704, n13707, n13708, n13709,
    n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
    n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13761, n13762, n13763, n13766,
    n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
    n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13788, n13789, n13791, n13792, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13818,
    n13819, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
    n13829, n13830, n13831, n13832, n13833, n13834, n13837, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13863, n13864, n13866, n13867, n13868, n13869, n13870,
    n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
    n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
    n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
    n13907, n13908, n13909, n13910;
  invx  g00000(.a(pi00), .O(n45));
  invx  g00001(.a(pi03), .O(n46));
  invx  g00002(.a(pi04), .O(n47));
  invx  g00003(.a(pi05), .O(n48));
  invx  g00004(.a(pi06), .O(n49));
  invx  g00005(.a(pi07), .O(n50));
  invx  g00006(.a(pi08), .O(n51));
  invx  g00007(.a(pi09), .O(n52));
  invx  g00008(.a(pi10), .O(n53));
  invx  g00009(.a(pi11), .O(n54));
  invx  g00010(.a(pi12), .O(n55));
  invx  g00011(.a(pi17), .O(n56));
  invx  g00012(.a(pi18), .O(n57));
  invx  g00013(.a(pi19), .O(n58));
  andx  g00014(.a(n58), .b(n57), .O(n59));
  andx  g00015(.a(n59), .b(n56), .O(n60));
  orx   g00016(.a(pi16), .b(pi15), .O(n61));
  invx  g00017(.a(n61), .O(n62));
  andx  g00018(.a(n62), .b(n60), .O(n63));
  invx  g00019(.a(pi13), .O(n64));
  invx  g00020(.a(pi14), .O(n65));
  andx  g00021(.a(n65), .b(n64), .O(n66));
  andx  g00022(.a(n66), .b(n63), .O(n67));
  andx  g00023(.a(n67), .b(n55), .O(n68));
  andx  g00024(.a(n68), .b(n54), .O(n69));
  andx  g00025(.a(n69), .b(n53), .O(n70));
  andx  g00026(.a(n70), .b(n52), .O(n71));
  andx  g00027(.a(n71), .b(n51), .O(n72));
  andx  g00028(.a(n72), .b(n50), .O(n73));
  andx  g00029(.a(n73), .b(n49), .O(n74));
  andx  g00030(.a(n74), .b(n48), .O(n75));
  andx  g00031(.a(n75), .b(n47), .O(n76));
  andx  g00032(.a(n76), .b(n46), .O(n77));
  invx  g00033(.a(pi01), .O(n78));
  invx  g00034(.a(pi02), .O(n79));
  andx  g00035(.a(n79), .b(n78), .O(n80));
  andx  g00036(.a(n80), .b(n77), .O(n81));
  andx  g00037(.a(n81), .b(n45), .O(n82));
  invx  g00038(.a(n82), .O(n83));
  invx  g00039(.a(n77), .O(n84));
  orx   g00040(.a(n84), .b(pi02), .O(n85));
  andx  g00041(.a(n73), .b(pi06), .O(n86));
  orx   g00042(.a(pi19), .b(pi18), .O(n87));
  orx   g00043(.a(n87), .b(pi17), .O(n88));
  orx   g00044(.a(n61), .b(n88), .O(po04));
  invx  g00045(.a(n66), .O(n90));
  orx   g00046(.a(n90), .b(po04), .O(n91));
  orx   g00047(.a(n91), .b(pi12), .O(n92));
  orx   g00048(.a(n92), .b(pi11), .O(n93));
  orx   g00049(.a(n93), .b(pi10), .O(n94));
  orx   g00050(.a(n94), .b(pi09), .O(n95));
  orx   g00051(.a(n95), .b(pi08), .O(n96));
  andx  g00052(.a(n70), .b(pi09), .O(n97));
  invx  g00053(.a(n97), .O(n98));
  andx  g00054(.a(n68), .b(pi11), .O(n99));
  invx  g00055(.a(n99), .O(n100));
  orx   g00056(.a(po04), .b(pi14), .O(n101));
  orx   g00057(.a(n101), .b(n67), .O(n102));
  andx  g00058(.a(n58), .b(pi18), .O(n103));
  orx   g00059(.a(n103), .b(n60), .O(n104));
  orx   g00060(.a(n88), .b(pi16), .O(n105));
  orx   g00061(.a(n105), .b(n63), .O(n106));
  andx  g00062(.a(n106), .b(n104), .O(n107));
  andx  g00063(.a(n107), .b(n102), .O(n108));
  andx  g00064(.a(n108), .b(n100), .O(n109));
  andx  g00065(.a(n109), .b(n98), .O(n110));
  andx  g00066(.a(n110), .b(n96), .O(n111));
  orx   g00067(.a(n111), .b(n86), .O(n112));
  orx   g00068(.a(n112), .b(n75), .O(n113));
  andx  g00069(.a(n76), .b(pi03), .O(n114));
  invx  g00070(.a(n114), .O(n115));
  andx  g00071(.a(n115), .b(n113), .O(n116));
  andx  g00072(.a(n116), .b(n85), .O(n117));
  orx   g00073(.a(n117), .b(n81), .O(n118));
  andx  g00074(.a(n118), .b(n83), .O(po00));
  invx  g00075(.a(n81), .O(n120));
  invx  g00076(.a(n75), .O(n121));
  andx  g00077(.a(n88), .b(n58), .O(n122));
  orx   g00078(.a(n122), .b(n63), .O(n123));
  andx  g00079(.a(n123), .b(n91), .O(n124));
  orx   g00080(.a(n124), .b(n69), .O(n125));
  andx  g00081(.a(n125), .b(n95), .O(n126));
  orx   g00082(.a(n126), .b(n73), .O(n127));
  andx  g00083(.a(n127), .b(n121), .O(n128));
  orx   g00084(.a(n128), .b(n77), .O(n129));
  andx  g00085(.a(n129), .b(n120), .O(po01));
  orx   g00086(.a(n63), .b(pi19), .O(n131));
  andx  g00087(.a(n131), .b(n93), .O(n132));
  orx   g00088(.a(n132), .b(n73), .O(n133));
  andx  g00089(.a(n133), .b(n84), .O(po02));
  orx   g00090(.a(n96), .b(pi07), .O(n135));
  andx  g00091(.a(n135), .b(n63), .O(po03));
  andx  g00092(.a(n71), .b(pi08), .O(n137));
  andx  g00093(.a(n137), .b(pi00), .O(n138));
  invx  g00094(.a(n138), .O(n139));
  andx  g00095(.a(n97), .b(pi01), .O(n140));
  invx  g00096(.a(n140), .O(n141));
  orx   g00097(.a(n93), .b(n53), .O(n142));
  invx  g00098(.a(n142), .O(n143));
  andx  g00099(.a(n143), .b(pi02), .O(n144));
  invx  g00100(.a(n144), .O(n145));
  andx  g00101(.a(n99), .b(pi03), .O(n146));
  invx  g00102(.a(n146), .O(n147));
  andx  g00103(.a(n63), .b(pi14), .O(n148));
  invx  g00104(.a(n148), .O(n149));
  orx   g00105(.a(n149), .b(n49), .O(n150));
  andx  g00106(.a(n67), .b(pi04), .O(n151));
  invx  g00107(.a(n105), .O(n152));
  andx  g00108(.a(n152), .b(po04), .O(n153));
  andx  g00109(.a(n153), .b(pi07), .O(n154));
  orx   g00110(.a(n154), .b(n151), .O(n155));
  invx  g00111(.a(n155), .O(n156));
  andx  g00112(.a(n156), .b(n150), .O(n157));
  invx  g00113(.a(n101), .O(n158));
  andx  g00114(.a(n158), .b(n91), .O(n159));
  andx  g00115(.a(n159), .b(pi05), .O(n160));
  andx  g00116(.a(n59), .b(pi17), .O(n161));
  andx  g00117(.a(n161), .b(pi09), .O(n162));
  invx  g00118(.a(pi16), .O(n163));
  orx   g00119(.a(n88), .b(n163), .O(n164));
  invx  g00120(.a(n164), .O(n165));
  andx  g00121(.a(n165), .b(pi08), .O(n166));
  andx  g00122(.a(pi19), .b(pi11), .O(n167));
  andx  g00123(.a(n103), .b(pi10), .O(n168));
  orx   g00124(.a(n168), .b(n167), .O(n169));
  orx   g00125(.a(n169), .b(n166), .O(n170));
  orx   g00126(.a(n170), .b(n162), .O(n171));
  orx   g00127(.a(n171), .b(n160), .O(n172));
  invx  g00128(.a(n172), .O(n173));
  andx  g00129(.a(n173), .b(n157), .O(n174));
  orx   g00130(.a(n174), .b(n68), .O(n175));
  andx  g00131(.a(n175), .b(n147), .O(n176));
  andx  g00132(.a(n176), .b(n145), .O(n177));
  andx  g00133(.a(n177), .b(n141), .O(n178));
  andx  g00134(.a(n178), .b(n139), .O(n179));
  orx   g00135(.a(n96), .b(n50), .O(n180));
  orx   g00136(.a(n180), .b(n45), .O(n181));
  invx  g00137(.a(n181), .O(n182));
  invx  g00138(.a(n137), .O(n183));
  orx   g00139(.a(n183), .b(n78), .O(n184));
  invx  g00140(.a(n184), .O(n185));
  orx   g00141(.a(n98), .b(n79), .O(n186));
  invx  g00142(.a(n186), .O(n187));
  orx   g00143(.a(n142), .b(n46), .O(n188));
  invx  g00144(.a(n188), .O(n189));
  orx   g00145(.a(n100), .b(n47), .O(n190));
  invx  g00146(.a(n190), .O(n191));
  andx  g00147(.a(n148), .b(pi07), .O(n192));
  andx  g00148(.a(n67), .b(pi05), .O(n193));
  andx  g00149(.a(n153), .b(pi08), .O(n194));
  orx   g00150(.a(n194), .b(n193), .O(n195));
  orx   g00151(.a(n195), .b(n192), .O(n196));
  andx  g00152(.a(n159), .b(pi06), .O(n197));
  invx  g00153(.a(n161), .O(n198));
  orx   g00154(.a(n198), .b(n53), .O(n199));
  invx  g00155(.a(n199), .O(n200));
  andx  g00156(.a(n165), .b(pi09), .O(n201));
  andx  g00157(.a(pi19), .b(pi12), .O(n202));
  andx  g00158(.a(n103), .b(pi11), .O(n203));
  orx   g00159(.a(n203), .b(n202), .O(n204));
  orx   g00160(.a(n204), .b(n201), .O(n205));
  orx   g00161(.a(n205), .b(n200), .O(n206));
  orx   g00162(.a(n206), .b(n197), .O(n207));
  orx   g00163(.a(n207), .b(n196), .O(n208));
  andx  g00164(.a(n208), .b(n92), .O(n209));
  orx   g00165(.a(n209), .b(n191), .O(n210));
  orx   g00166(.a(n210), .b(n189), .O(n211));
  orx   g00167(.a(n211), .b(n187), .O(n212));
  orx   g00168(.a(n212), .b(n185), .O(n213));
  orx   g00169(.a(n213), .b(n182), .O(n214));
  invx  g00170(.a(n214), .O(n215));
  andx  g00171(.a(n215), .b(n179), .O(n216));
  invx  g00172(.a(n86), .O(n217));
  orx   g00173(.a(n217), .b(n45), .O(n218));
  orx   g00174(.a(n180), .b(n78), .O(n219));
  orx   g00175(.a(n183), .b(n79), .O(n220));
  orx   g00176(.a(n98), .b(n46), .O(n221));
  orx   g00177(.a(n149), .b(n51), .O(n222));
  andx  g00178(.a(n67), .b(pi06), .O(n223));
  andx  g00179(.a(n153), .b(pi09), .O(n224));
  orx   g00180(.a(n224), .b(n223), .O(n225));
  invx  g00181(.a(n225), .O(n226));
  andx  g00182(.a(n226), .b(n222), .O(n227));
  andx  g00183(.a(n159), .b(pi07), .O(n228));
  andx  g00184(.a(n161), .b(pi11), .O(n229));
  andx  g00185(.a(n165), .b(pi10), .O(n230));
  andx  g00186(.a(pi19), .b(pi13), .O(n231));
  andx  g00187(.a(n103), .b(pi12), .O(n232));
  orx   g00188(.a(n232), .b(n231), .O(n233));
  orx   g00189(.a(n233), .b(n230), .O(n234));
  orx   g00190(.a(n234), .b(n229), .O(n235));
  orx   g00191(.a(n235), .b(n228), .O(n236));
  invx  g00192(.a(n236), .O(n237));
  andx  g00193(.a(n237), .b(n227), .O(n238));
  orx   g00194(.a(n238), .b(n68), .O(n239));
  orx   g00195(.a(n100), .b(n48), .O(n240));
  andx  g00196(.a(n143), .b(pi04), .O(n241));
  invx  g00197(.a(n241), .O(n242));
  andx  g00198(.a(n242), .b(n240), .O(n243));
  andx  g00199(.a(n243), .b(n239), .O(n244));
  andx  g00200(.a(n244), .b(n221), .O(n245));
  andx  g00201(.a(n245), .b(n220), .O(n246));
  andx  g00202(.a(n246), .b(n219), .O(n247));
  andx  g00203(.a(n247), .b(n218), .O(n248));
  andx  g00204(.a(n248), .b(n216), .O(n249));
  invx  g00205(.a(n179), .O(n250));
  orx   g00206(.a(n214), .b(n250), .O(n251));
  invx  g00207(.a(n248), .O(n252));
  andx  g00208(.a(n252), .b(n251), .O(n253));
  orx   g00209(.a(n253), .b(n249), .O(n254));
  invx  g00210(.a(n254), .O(n255));
  andx  g00211(.a(n77), .b(pi00), .O(n256));
  andx  g00212(.a(n75), .b(pi04), .O(n257));
  orx   g00213(.a(n257), .b(n256), .O(n258));
  andx  g00214(.a(n258), .b(pi02), .O(n259));
  andx  g00215(.a(n114), .b(pi01), .O(n260));
  orx   g00216(.a(n217), .b(n47), .O(n261));
  invx  g00217(.a(n261), .O(n262));
  orx   g00218(.a(n183), .b(n49), .O(n263));
  orx   g00219(.a(n98), .b(n50), .O(n264));
  orx   g00220(.a(n149), .b(n55), .O(n265));
  andx  g00221(.a(n67), .b(pi10), .O(n266));
  andx  g00222(.a(n153), .b(pi13), .O(n267));
  orx   g00223(.a(n267), .b(n266), .O(n268));
  invx  g00224(.a(n268), .O(n269));
  andx  g00225(.a(n269), .b(n265), .O(n270));
  andx  g00226(.a(n159), .b(pi11), .O(n271));
  andx  g00227(.a(n161), .b(pi15), .O(n272));
  andx  g00228(.a(n165), .b(pi14), .O(n273));
  andx  g00229(.a(pi19), .b(pi17), .O(n274));
  andx  g00230(.a(n103), .b(pi16), .O(n275));
  orx   g00231(.a(n275), .b(n274), .O(n276));
  orx   g00232(.a(n276), .b(n273), .O(n277));
  orx   g00233(.a(n277), .b(n272), .O(n278));
  orx   g00234(.a(n278), .b(n271), .O(n279));
  invx  g00235(.a(n279), .O(n280));
  andx  g00236(.a(n280), .b(n270), .O(n281));
  orx   g00237(.a(n281), .b(n68), .O(n282));
  andx  g00238(.a(n143), .b(pi08), .O(n283));
  invx  g00239(.a(n283), .O(n284));
  orx   g00240(.a(n100), .b(n52), .O(n285));
  andx  g00241(.a(n285), .b(n284), .O(n286));
  andx  g00242(.a(n286), .b(n282), .O(n287));
  andx  g00243(.a(n287), .b(n264), .O(n288));
  andx  g00244(.a(n288), .b(n263), .O(n289));
  invx  g00245(.a(n289), .O(n290));
  invx  g00246(.a(n180), .O(n291));
  andx  g00247(.a(n291), .b(pi05), .O(n292));
  andx  g00248(.a(n74), .b(pi03), .O(n293));
  orx   g00249(.a(n293), .b(n292), .O(n294));
  orx   g00250(.a(n294), .b(n290), .O(n295));
  orx   g00251(.a(n295), .b(n262), .O(n296));
  andx  g00252(.a(n296), .b(n121), .O(n297));
  orx   g00253(.a(n297), .b(n260), .O(n298));
  orx   g00254(.a(n298), .b(n259), .O(n299));
  andx  g00255(.a(n299), .b(n250), .O(n300));
  andx  g00256(.a(n114), .b(pi00), .O(n301));
  andx  g00257(.a(n257), .b(pi01), .O(n302));
  andx  g00258(.a(n86), .b(pi03), .O(n303));
  andx  g00259(.a(n137), .b(pi05), .O(n304));
  andx  g00260(.a(n97), .b(pi06), .O(n305));
  andx  g00261(.a(n148), .b(pi11), .O(n306));
  andx  g00262(.a(n67), .b(pi09), .O(n307));
  andx  g00263(.a(n153), .b(pi12), .O(n308));
  orx   g00264(.a(n308), .b(n307), .O(n309));
  orx   g00265(.a(n309), .b(n306), .O(n310));
  andx  g00266(.a(n159), .b(pi10), .O(n311));
  orx   g00267(.a(n198), .b(n65), .O(n312));
  invx  g00268(.a(n312), .O(n313));
  andx  g00269(.a(n165), .b(pi13), .O(n314));
  andx  g00270(.a(pi19), .b(pi16), .O(n315));
  andx  g00271(.a(n103), .b(pi15), .O(n316));
  orx   g00272(.a(n316), .b(n315), .O(n317));
  orx   g00273(.a(n317), .b(n314), .O(n318));
  orx   g00274(.a(n318), .b(n313), .O(n319));
  orx   g00275(.a(n319), .b(n311), .O(n320));
  orx   g00276(.a(n320), .b(n310), .O(n321));
  andx  g00277(.a(n321), .b(n92), .O(n322));
  andx  g00278(.a(n143), .b(pi07), .O(n323));
  andx  g00279(.a(n99), .b(pi08), .O(n324));
  orx   g00280(.a(n324), .b(n323), .O(n325));
  orx   g00281(.a(n325), .b(n322), .O(n326));
  orx   g00282(.a(n326), .b(n305), .O(n327));
  orx   g00283(.a(n327), .b(n304), .O(n328));
  andx  g00284(.a(n291), .b(pi04), .O(n329));
  orx   g00285(.a(n135), .b(pi06), .O(n330));
  orx   g00286(.a(n330), .b(n79), .O(n331));
  invx  g00287(.a(n331), .O(n332));
  orx   g00288(.a(n332), .b(n329), .O(n333));
  orx   g00289(.a(n333), .b(n328), .O(n334));
  orx   g00290(.a(n334), .b(n303), .O(n335));
  andx  g00291(.a(n335), .b(n121), .O(n336));
  orx   g00292(.a(n336), .b(n302), .O(n337));
  orx   g00293(.a(n337), .b(n301), .O(n338));
  andx  g00294(.a(n338), .b(n250), .O(n339));
  andx  g00295(.a(n86), .b(pi02), .O(n340));
  andx  g00296(.a(n137), .b(pi04), .O(n341));
  andx  g00297(.a(n97), .b(pi05), .O(n342));
  andx  g00298(.a(n148), .b(pi10), .O(n343));
  orx   g00299(.a(n91), .b(n51), .O(n344));
  invx  g00300(.a(n344), .O(n345));
  andx  g00301(.a(n153), .b(pi11), .O(n346));
  orx   g00302(.a(n346), .b(n345), .O(n347));
  orx   g00303(.a(n347), .b(n343), .O(n348));
  andx  g00304(.a(n159), .b(pi09), .O(n349));
  andx  g00305(.a(n161), .b(pi13), .O(n350));
  orx   g00306(.a(n164), .b(n55), .O(n351));
  invx  g00307(.a(n351), .O(n352));
  andx  g00308(.a(pi19), .b(pi15), .O(n353));
  andx  g00309(.a(n103), .b(pi14), .O(n354));
  orx   g00310(.a(n354), .b(n353), .O(n355));
  orx   g00311(.a(n355), .b(n352), .O(n356));
  orx   g00312(.a(n356), .b(n350), .O(n357));
  orx   g00313(.a(n357), .b(n349), .O(n358));
  orx   g00314(.a(n358), .b(n348), .O(n359));
  andx  g00315(.a(n359), .b(n92), .O(n360));
  orx   g00316(.a(n142), .b(n49), .O(n361));
  invx  g00317(.a(n361), .O(n362));
  andx  g00318(.a(n99), .b(pi07), .O(n363));
  orx   g00319(.a(n363), .b(n362), .O(n364));
  orx   g00320(.a(n364), .b(n360), .O(n365));
  orx   g00321(.a(n365), .b(n342), .O(n366));
  orx   g00322(.a(n366), .b(n341), .O(n367));
  orx   g00323(.a(n180), .b(n46), .O(n368));
  invx  g00324(.a(n368), .O(n369));
  andx  g00325(.a(n74), .b(pi01), .O(n370));
  orx   g00326(.a(n370), .b(n369), .O(n371));
  orx   g00327(.a(n371), .b(n367), .O(n372));
  orx   g00328(.a(n372), .b(n340), .O(n373));
  andx  g00329(.a(n373), .b(n121), .O(n374));
  andx  g00330(.a(n257), .b(pi00), .O(n375));
  orx   g00331(.a(n375), .b(n374), .O(n376));
  andx  g00332(.a(n214), .b(n250), .O(n377));
  orx   g00333(.a(n377), .b(n216), .O(n378));
  invx  g00334(.a(n378), .O(n379));
  andx  g00335(.a(n379), .b(n376), .O(n380));
  invx  g00336(.a(n380), .O(n381));
  andx  g00337(.a(n97), .b(pi00), .O(n382));
  andx  g00338(.a(n143), .b(pi01), .O(n383));
  andx  g00339(.a(n148), .b(pi05), .O(n384));
  andx  g00340(.a(n153), .b(pi06), .O(n385));
  andx  g00341(.a(n67), .b(pi03), .O(n386));
  orx   g00342(.a(n386), .b(n385), .O(n387));
  orx   g00343(.a(n387), .b(n384), .O(n388));
  andx  g00344(.a(n159), .b(pi04), .O(n389));
  andx  g00345(.a(n165), .b(pi07), .O(n390));
  andx  g00346(.a(n161), .b(pi08), .O(n391));
  andx  g00347(.a(n103), .b(pi09), .O(n392));
  andx  g00348(.a(pi19), .b(pi10), .O(n393));
  orx   g00349(.a(n393), .b(n392), .O(n394));
  orx   g00350(.a(n394), .b(n391), .O(n395));
  orx   g00351(.a(n395), .b(n390), .O(n396));
  orx   g00352(.a(n396), .b(n389), .O(n397));
  orx   g00353(.a(n397), .b(n388), .O(n398));
  andx  g00354(.a(n398), .b(n92), .O(n399));
  andx  g00355(.a(n99), .b(pi02), .O(n400));
  orx   g00356(.a(n400), .b(n399), .O(n401));
  orx   g00357(.a(n401), .b(n383), .O(n402));
  orx   g00358(.a(n402), .b(n382), .O(n403));
  invx  g00359(.a(n403), .O(n404));
  orx   g00360(.a(n252), .b(n251), .O(n405));
  andx  g00361(.a(n86), .b(pi01), .O(n406));
  andx  g00362(.a(n137), .b(pi03), .O(n407));
  andx  g00363(.a(n97), .b(pi04), .O(n408));
  andx  g00364(.a(n148), .b(pi09), .O(n409));
  andx  g00365(.a(n67), .b(pi07), .O(n410));
  andx  g00366(.a(n153), .b(pi10), .O(n411));
  orx   g00367(.a(n411), .b(n410), .O(n412));
  orx   g00368(.a(n412), .b(n409), .O(n413));
  andx  g00369(.a(n159), .b(pi08), .O(n414));
  orx   g00370(.a(n198), .b(n55), .O(n415));
  invx  g00371(.a(n415), .O(n416));
  andx  g00372(.a(n165), .b(pi11), .O(n417));
  andx  g00373(.a(pi19), .b(pi14), .O(n418));
  andx  g00374(.a(n103), .b(pi13), .O(n419));
  orx   g00375(.a(n419), .b(n418), .O(n420));
  orx   g00376(.a(n420), .b(n417), .O(n421));
  orx   g00377(.a(n421), .b(n416), .O(n422));
  orx   g00378(.a(n422), .b(n414), .O(n423));
  orx   g00379(.a(n423), .b(n413), .O(n424));
  andx  g00380(.a(n424), .b(n92), .O(n425));
  andx  g00381(.a(n143), .b(pi05), .O(n426));
  andx  g00382(.a(n99), .b(pi06), .O(n427));
  orx   g00383(.a(n427), .b(n426), .O(n428));
  orx   g00384(.a(n428), .b(n425), .O(n429));
  orx   g00385(.a(n429), .b(n408), .O(n430));
  orx   g00386(.a(n430), .b(n407), .O(n431));
  andx  g00387(.a(n291), .b(pi02), .O(n432));
  orx   g00388(.a(n330), .b(n45), .O(n433));
  invx  g00389(.a(n433), .O(n434));
  orx   g00390(.a(n434), .b(n432), .O(n435));
  orx   g00391(.a(n435), .b(n431), .O(n436));
  orx   g00392(.a(n436), .b(n406), .O(n437));
  andx  g00393(.a(n437), .b(n121), .O(n438));
  orx   g00394(.a(n438), .b(n405), .O(n439));
  andx  g00395(.a(n439), .b(n376), .O(n440));
  invx  g00396(.a(n340), .O(n441));
  invx  g00397(.a(n341), .O(n442));
  invx  g00398(.a(n342), .O(n443));
  invx  g00399(.a(n343), .O(n444));
  orx   g00400(.a(n106), .b(n54), .O(n445));
  andx  g00401(.a(n445), .b(n344), .O(n446));
  andx  g00402(.a(n446), .b(n444), .O(n447));
  orx   g00403(.a(n102), .b(n52), .O(n448));
  invx  g00404(.a(n350), .O(n449));
  invx  g00405(.a(n355), .O(n450));
  andx  g00406(.a(n450), .b(n351), .O(n451));
  andx  g00407(.a(n451), .b(n449), .O(n452));
  andx  g00408(.a(n452), .b(n448), .O(n453));
  andx  g00409(.a(n453), .b(n447), .O(n454));
  orx   g00410(.a(n454), .b(n68), .O(n455));
  invx  g00411(.a(n363), .O(n456));
  andx  g00412(.a(n456), .b(n361), .O(n457));
  andx  g00413(.a(n457), .b(n455), .O(n458));
  andx  g00414(.a(n458), .b(n443), .O(n459));
  andx  g00415(.a(n459), .b(n442), .O(n460));
  orx   g00416(.a(n330), .b(n78), .O(n461));
  andx  g00417(.a(n461), .b(n368), .O(n462));
  andx  g00418(.a(n462), .b(n460), .O(n463));
  andx  g00419(.a(n463), .b(n441), .O(n464));
  orx   g00420(.a(n464), .b(n75), .O(n465));
  invx  g00421(.a(n375), .O(n466));
  andx  g00422(.a(n466), .b(n465), .O(n467));
  invx  g00423(.a(n406), .O(n468));
  invx  g00424(.a(n431), .O(n469));
  invx  g00425(.a(n432), .O(n470));
  andx  g00426(.a(n433), .b(n470), .O(n471));
  andx  g00427(.a(n471), .b(n469), .O(n472));
  andx  g00428(.a(n472), .b(n468), .O(n473));
  orx   g00429(.a(n473), .b(n75), .O(n474));
  andx  g00430(.a(n474), .b(n467), .O(n475));
  andx  g00431(.a(n475), .b(n249), .O(n476));
  orx   g00432(.a(n476), .b(n440), .O(n477));
  orx   g00433(.a(n477), .b(n404), .O(n478));
  andx  g00434(.a(n474), .b(n249), .O(n479));
  andx  g00435(.a(n438), .b(n405), .O(n480));
  orx   g00436(.a(n480), .b(n479), .O(n481));
  orx   g00437(.a(n481), .b(n179), .O(n482));
  invx  g00438(.a(n482), .O(n483));
  andx  g00439(.a(n483), .b(n478), .O(n484));
  orx   g00440(.a(n479), .b(n467), .O(n485));
  orx   g00441(.a(n438), .b(n376), .O(n486));
  orx   g00442(.a(n486), .b(n405), .O(n487));
  andx  g00443(.a(n487), .b(n485), .O(n488));
  andx  g00444(.a(n488), .b(n403), .O(n489));
  andx  g00445(.a(n482), .b(n489), .O(n490));
  orx   g00446(.a(n490), .b(n484), .O(n491));
  andx  g00447(.a(n255), .b(n214), .O(n492));
  orx   g00448(.a(n492), .b(n491), .O(n493));
  andx  g00449(.a(n492), .b(n491), .O(n494));
  invx  g00450(.a(n494), .O(n495));
  andx  g00451(.a(n495), .b(n493), .O(n496));
  orx   g00452(.a(n254), .b(n179), .O(n497));
  invx  g00453(.a(n497), .O(n498));
  invx  g00454(.a(n481), .O(n499));
  andx  g00455(.a(n499), .b(n403), .O(n500));
  orx   g00456(.a(n500), .b(n498), .O(n501));
  andx  g00457(.a(n500), .b(n498), .O(n502));
  invx  g00458(.a(n502), .O(n503));
  andx  g00459(.a(n503), .b(n501), .O(n504));
  andx  g00460(.a(n403), .b(n379), .O(n505));
  andx  g00461(.a(n505), .b(n498), .O(n506));
  andx  g00462(.a(n506), .b(n504), .O(n507));
  andx  g00463(.a(n214), .b(n179), .O(n508));
  andx  g00464(.a(n508), .b(n504), .O(n509));
  orx   g00465(.a(n509), .b(n507), .O(n510));
  andx  g00466(.a(n510), .b(n496), .O(n511));
  invx  g00467(.a(n511), .O(n512));
  andx  g00468(.a(n379), .b(n252), .O(n513));
  invx  g00469(.a(n513), .O(n514));
  invx  g00470(.a(n493), .O(n515));
  orx   g00471(.a(n494), .b(n515), .O(n516));
  invx  g00472(.a(n501), .O(n517));
  orx   g00473(.a(n502), .b(n517), .O(n518));
  invx  g00474(.a(n506), .O(n519));
  orx   g00475(.a(n519), .b(n518), .O(n520));
  invx  g00476(.a(n508), .O(n521));
  orx   g00477(.a(n521), .b(n518), .O(n522));
  andx  g00478(.a(n522), .b(n520), .O(n523));
  andx  g00479(.a(n523), .b(n516), .O(n524));
  orx   g00480(.a(n524), .b(n514), .O(n525));
  andx  g00481(.a(n525), .b(n512), .O(n526));
  andx  g00482(.a(n502), .b(n214), .O(n527));
  invx  g00483(.a(n527), .O(n528));
  invx  g00484(.a(n491), .O(n529));
  invx  g00485(.a(n492), .O(n530));
  andx  g00486(.a(n503), .b(n530), .O(n531));
  orx   g00487(.a(n531), .b(n529), .O(n532));
  andx  g00488(.a(n532), .b(n528), .O(n533));
  invx  g00489(.a(n533), .O(n534));
  andx  g00490(.a(n483), .b(n489), .O(n535));
  andx  g00491(.a(n499), .b(n214), .O(n536));
  orx   g00492(.a(n536), .b(n535), .O(n537));
  andx  g00493(.a(n535), .b(n214), .O(n538));
  invx  g00494(.a(n538), .O(n539));
  andx  g00495(.a(n539), .b(n537), .O(n540));
  invx  g00496(.a(n301), .O(n541));
  invx  g00497(.a(n302), .O(n542));
  invx  g00498(.a(n303), .O(n543));
  invx  g00499(.a(n328), .O(n544));
  invx  g00500(.a(n329), .O(n545));
  andx  g00501(.a(n331), .b(n545), .O(n546));
  andx  g00502(.a(n546), .b(n544), .O(n547));
  andx  g00503(.a(n547), .b(n543), .O(n548));
  orx   g00504(.a(n548), .b(n75), .O(n549));
  andx  g00505(.a(n549), .b(n542), .O(n550));
  andx  g00506(.a(n550), .b(n541), .O(n551));
  orx   g00507(.a(n476), .b(n551), .O(n552));
  orx   g00508(.a(n487), .b(n338), .O(n553));
  andx  g00509(.a(n553), .b(n552), .O(n554));
  andx  g00510(.a(n554), .b(n403), .O(n555));
  orx   g00511(.a(n477), .b(n179), .O(n556));
  orx   g00512(.a(n556), .b(n555), .O(n557));
  andx  g00513(.a(n487), .b(n338), .O(n558));
  andx  g00514(.a(n476), .b(n551), .O(n559));
  orx   g00515(.a(n559), .b(n558), .O(n560));
  orx   g00516(.a(n560), .b(n404), .O(n561));
  andx  g00517(.a(n488), .b(n250), .O(n562));
  orx   g00518(.a(n562), .b(n561), .O(n563));
  andx  g00519(.a(n563), .b(n557), .O(n564));
  orx   g00520(.a(n564), .b(n540), .O(n565));
  invx  g00521(.a(n565), .O(n566));
  andx  g00522(.a(n564), .b(n540), .O(n567));
  orx   g00523(.a(n567), .b(n566), .O(n568));
  andx  g00524(.a(n568), .b(n534), .O(n569));
  invx  g00525(.a(n567), .O(n570));
  andx  g00526(.a(n570), .b(n565), .O(n571));
  andx  g00527(.a(n571), .b(n533), .O(n572));
  orx   g00528(.a(n572), .b(n569), .O(n573));
  andx  g00529(.a(n573), .b(n526), .O(n574));
  invx  g00530(.a(n574), .O(n575));
  orx   g00531(.a(n510), .b(n496), .O(n576));
  andx  g00532(.a(n576), .b(n513), .O(n577));
  orx   g00533(.a(n577), .b(n511), .O(n578));
  andx  g00534(.a(n438), .b(n379), .O(n579));
  orx   g00535(.a(n579), .b(n578), .O(n580));
  orx   g00536(.a(n571), .b(n533), .O(n581));
  orx   g00537(.a(n568), .b(n534), .O(n582));
  andx  g00538(.a(n582), .b(n581), .O(n583));
  orx   g00539(.a(n579), .b(n583), .O(n584));
  andx  g00540(.a(n584), .b(n580), .O(n585));
  andx  g00541(.a(n585), .b(n575), .O(n586));
  orx   g00542(.a(n586), .b(n381), .O(n587));
  invx  g00543(.a(n579), .O(n588));
  andx  g00544(.a(n588), .b(n526), .O(n589));
  andx  g00545(.a(n588), .b(n573), .O(n590));
  orx   g00546(.a(n590), .b(n589), .O(n591));
  orx   g00547(.a(n591), .b(n574), .O(n592));
  orx   g00548(.a(n592), .b(n380), .O(n593));
  andx  g00549(.a(n593), .b(n587), .O(n594));
  invx  g00550(.a(n259), .O(n595));
  invx  g00551(.a(n260), .O(n596));
  invx  g00552(.a(n294), .O(n597));
  andx  g00553(.a(n597), .b(n289), .O(n598));
  andx  g00554(.a(n598), .b(n261), .O(n599));
  orx   g00555(.a(n599), .b(n75), .O(n600));
  andx  g00556(.a(n600), .b(n596), .O(n601));
  andx  g00557(.a(n601), .b(n595), .O(n602));
  orx   g00558(.a(n559), .b(n602), .O(n603));
  orx   g00559(.a(n553), .b(n299), .O(n604));
  andx  g00560(.a(n604), .b(n603), .O(n605));
  andx  g00561(.a(n605), .b(n403), .O(n606));
  orx   g00562(.a(n560), .b(n179), .O(n607));
  orx   g00563(.a(n607), .b(n606), .O(n608));
  andx  g00564(.a(n553), .b(n299), .O(n609));
  andx  g00565(.a(n559), .b(n602), .O(n610));
  orx   g00566(.a(n610), .b(n609), .O(n611));
  orx   g00567(.a(n611), .b(n404), .O(n612));
  andx  g00568(.a(n554), .b(n250), .O(n613));
  orx   g00569(.a(n613), .b(n612), .O(n614));
  andx  g00570(.a(n614), .b(n608), .O(n615));
  andx  g00571(.a(n562), .b(n555), .O(n616));
  andx  g00572(.a(n488), .b(n214), .O(n617));
  invx  g00573(.a(n617), .O(n618));
  orx   g00574(.a(n618), .b(n616), .O(n619));
  orx   g00575(.a(n556), .b(n561), .O(n620));
  orx   g00576(.a(n617), .b(n620), .O(n621));
  andx  g00577(.a(n621), .b(n619), .O(n622));
  andx  g00578(.a(n622), .b(n615), .O(n623));
  andx  g00579(.a(n613), .b(n612), .O(n624));
  andx  g00580(.a(n607), .b(n606), .O(n625));
  orx   g00581(.a(n625), .b(n624), .O(n626));
  andx  g00582(.a(n617), .b(n620), .O(n627));
  andx  g00583(.a(n618), .b(n616), .O(n628));
  orx   g00584(.a(n628), .b(n627), .O(n629));
  andx  g00585(.a(n629), .b(n626), .O(n630));
  orx   g00586(.a(n630), .b(n623), .O(n631));
  andx  g00587(.a(n499), .b(n252), .O(n632));
  invx  g00588(.a(n632), .O(n633));
  andx  g00589(.a(n562), .b(n561), .O(n634));
  andx  g00590(.a(n556), .b(n555), .O(n635));
  orx   g00591(.a(n635), .b(n634), .O(n636));
  andx  g00592(.a(n636), .b(n537), .O(n637));
  orx   g00593(.a(n637), .b(n538), .O(n638));
  andx  g00594(.a(n638), .b(n633), .O(n639));
  orx   g00595(.a(n482), .b(n478), .O(n640));
  invx  g00596(.a(n536), .O(n641));
  andx  g00597(.a(n641), .b(n640), .O(n642));
  orx   g00598(.a(n564), .b(n642), .O(n643));
  andx  g00599(.a(n643), .b(n539), .O(n644));
  andx  g00600(.a(n644), .b(n632), .O(n645));
  orx   g00601(.a(n645), .b(n639), .O(n646));
  andx  g00602(.a(n646), .b(n631), .O(n647));
  orx   g00603(.a(n629), .b(n626), .O(n648));
  orx   g00604(.a(n622), .b(n615), .O(n649));
  andx  g00605(.a(n649), .b(n648), .O(n650));
  orx   g00606(.a(n644), .b(n632), .O(n651));
  orx   g00607(.a(n638), .b(n633), .O(n652));
  andx  g00608(.a(n652), .b(n651), .O(n653));
  andx  g00609(.a(n653), .b(n650), .O(n654));
  orx   g00610(.a(n654), .b(n647), .O(n655));
  andx  g00611(.a(n438), .b(n255), .O(n656));
  invx  g00612(.a(n656), .O(n657));
  andx  g00613(.a(n252), .b(n216), .O(n658));
  invx  g00614(.a(n658), .O(n659));
  andx  g00615(.a(n659), .b(n533), .O(n660));
  orx   g00616(.a(n660), .b(n571), .O(n661));
  andx  g00617(.a(n661), .b(n657), .O(n662));
  invx  g00618(.a(n660), .O(n663));
  andx  g00619(.a(n663), .b(n568), .O(n664));
  andx  g00620(.a(n664), .b(n656), .O(n665));
  orx   g00621(.a(n665), .b(n662), .O(n666));
  andx  g00622(.a(n666), .b(n655), .O(n667));
  orx   g00623(.a(n653), .b(n650), .O(n668));
  orx   g00624(.a(n646), .b(n631), .O(n669));
  andx  g00625(.a(n669), .b(n668), .O(n670));
  orx   g00626(.a(n664), .b(n656), .O(n671));
  orx   g00627(.a(n661), .b(n657), .O(n672));
  andx  g00628(.a(n672), .b(n671), .O(n673));
  andx  g00629(.a(n673), .b(n670), .O(n674));
  orx   g00630(.a(n674), .b(n667), .O(n675));
  andx  g00631(.a(n675), .b(n594), .O(n676));
  andx  g00632(.a(n592), .b(n380), .O(n677));
  andx  g00633(.a(n586), .b(n381), .O(n678));
  orx   g00634(.a(n678), .b(n677), .O(n679));
  orx   g00635(.a(n673), .b(n670), .O(n680));
  orx   g00636(.a(n666), .b(n655), .O(n681));
  andx  g00637(.a(n681), .b(n680), .O(n682));
  andx  g00638(.a(n682), .b(n679), .O(n683));
  orx   g00639(.a(n683), .b(n676), .O(n684));
  orx   g00640(.a(n684), .b(n339), .O(n685));
  orx   g00641(.a(n588), .b(n526), .O(n686));
  andx  g00642(.a(n686), .b(n580), .O(n687));
  andx  g00643(.a(n583), .b(n687), .O(n691));
  andx  g00644(.a(n579), .b(n578), .O(n692));
  orx   g00645(.a(n692), .b(n589), .O(n693));
  andx  g00646(.a(n573), .b(n693), .O(n695));
  orx   g00647(.a(n695), .b(n691), .O(n696));
  andx  g00648(.a(n696), .b(n467), .O(n697));
  invx  g00649(.a(n697), .O(n698));
  orx   g00650(.a(n573), .b(n693), .O(n699));
  orx   g00651(.a(n583), .b(n687), .O(n700));
  andx  g00652(.a(n700), .b(n699), .O(n701));
  andx  g00653(.a(n701), .b(n376), .O(n702));
  andx  g00654(.a(n514), .b(n523), .O(n703));
  invx  g00655(.a(n703), .O(n704));
  andx  g00656(.a(n704), .b(n516), .O(n705));
  andx  g00657(.a(n703), .b(n496), .O(n706));
  orx   g00658(.a(n706), .b(n705), .O(n707));
  orx   g00659(.a(n707), .b(n702), .O(n708));
  orx   g00660(.a(n701), .b(n438), .O(n709));
  andx  g00661(.a(n486), .b(n250), .O(n710));
  andx  g00662(.a(n710), .b(n709), .O(n711));
  andx  g00663(.a(n711), .b(n708), .O(n712));
  invx  g00664(.a(n707), .O(n713));
  andx  g00665(.a(n713), .b(n474), .O(n714));
  invx  g00666(.a(n714), .O(n715));
  andx  g00667(.a(n252), .b(n250), .O(n716));
  andx  g00668(.a(n378), .b(n255), .O(n718));
  orx   g00669(.a(n718), .b(n513), .O(n719));
  andx  g00670(.a(n403), .b(n250), .O(n720));
  andx  g00671(.a(n720), .b(n719), .O(n721));
  andx  g00672(.a(n721), .b(n716), .O(n722));
  orx   g00673(.a(n722), .b(n504), .O(n723));
  orx   g00674(.a(n721), .b(n716), .O(n724));
  andx  g00675(.a(n724), .b(n723), .O(n725));
  andx  g00676(.a(n725), .b(n715), .O(n726));
  orx   g00677(.a(n726), .b(n712), .O(n727));
  andx  g00678(.a(n727), .b(n698), .O(n728));
  andx  g00679(.a(n728), .b(n685), .O(n729));
  andx  g00680(.a(n684), .b(n339), .O(n730));
  orx   g00681(.a(n730), .b(n729), .O(n731));
  andx  g00682(.a(n731), .b(n300), .O(n732));
  invx  g00683(.a(n300), .O(n733));
  invx  g00684(.a(n339), .O(n734));
  orx   g00685(.a(n682), .b(n679), .O(n735));
  orx   g00686(.a(n675), .b(n594), .O(n736));
  andx  g00687(.a(n736), .b(n735), .O(n737));
  andx  g00688(.a(n737), .b(n734), .O(n738));
  orx   g00689(.a(n696), .b(n467), .O(n739));
  andx  g00690(.a(n713), .b(n739), .O(n740));
  andx  g00691(.a(n696), .b(n474), .O(n741));
  invx  g00692(.a(n710), .O(n742));
  orx   g00693(.a(n742), .b(n741), .O(n743));
  orx   g00694(.a(n743), .b(n740), .O(n744));
  invx  g00695(.a(n726), .O(n745));
  andx  g00696(.a(n745), .b(n744), .O(n746));
  orx   g00697(.a(n746), .b(n697), .O(n747));
  orx   g00698(.a(n747), .b(n738), .O(n748));
  invx  g00699(.a(n730), .O(n749));
  andx  g00700(.a(n749), .b(n748), .O(n750));
  andx  g00701(.a(n750), .b(n733), .O(n751));
  orx   g00702(.a(n751), .b(n732), .O(n752));
  andx  g00703(.a(n376), .b(n255), .O(n753));
  orx   g00704(.a(n664), .b(n655), .O(n754));
  andx  g00705(.a(n664), .b(n655), .O(n755));
  orx   g00706(.a(n755), .b(n656), .O(n756));
  andx  g00707(.a(n756), .b(n754), .O(n757));
  andx  g00708(.a(n757), .b(n753), .O(n758));
  invx  g00709(.a(n753), .O(n759));
  andx  g00710(.a(n661), .b(n670), .O(n760));
  orx   g00711(.a(n661), .b(n670), .O(n761));
  andx  g00712(.a(n761), .b(n657), .O(n762));
  orx   g00713(.a(n762), .b(n760), .O(n763));
  andx  g00714(.a(n763), .b(n759), .O(n764));
  orx   g00715(.a(n764), .b(n758), .O(n765));
  andx  g00716(.a(n438), .b(n249), .O(n766));
  andx  g00717(.a(n650), .b(n632), .O(n770));
  andx  g00718(.a(n650), .b(n638), .O(n771));
  andx  g00719(.a(n638), .b(n632), .O(n772));
  orx   g00720(.a(n772), .b(n771), .O(n773));
  orx   g00721(.a(n773), .b(n770), .O(n774));
  orx   g00722(.a(n774), .b(n766), .O(n775));
  invx  g00723(.a(n775), .O(n776));
  andx  g00724(.a(n605), .b(n250), .O(n777));
  andx  g00725(.a(n86), .b(pi05), .O(n778));
  invx  g00726(.a(n778), .O(n779));
  andx  g00727(.a(n137), .b(pi07), .O(n780));
  invx  g00728(.a(n780), .O(n781));
  andx  g00729(.a(n97), .b(pi08), .O(n782));
  invx  g00730(.a(n782), .O(n783));
  andx  g00731(.a(n143), .b(pi09), .O(n784));
  invx  g00732(.a(n784), .O(n785));
  andx  g00733(.a(n148), .b(pi13), .O(n786));
  invx  g00734(.a(n786), .O(n787));
  andx  g00735(.a(n153), .b(pi14), .O(n788));
  invx  g00736(.a(n788), .O(n789));
  orx   g00737(.a(n91), .b(n54), .O(n790));
  andx  g00738(.a(n790), .b(n789), .O(n791));
  andx  g00739(.a(n791), .b(n787), .O(n792));
  andx  g00740(.a(n159), .b(pi12), .O(n793));
  andx  g00741(.a(n165), .b(pi15), .O(n794));
  andx  g00742(.a(n161), .b(pi16), .O(n795));
  andx  g00743(.a(n103), .b(pi17), .O(n796));
  andx  g00744(.a(pi19), .b(pi18), .O(n797));
  orx   g00745(.a(n797), .b(n796), .O(n798));
  orx   g00746(.a(n798), .b(n795), .O(n799));
  orx   g00747(.a(n799), .b(n794), .O(n800));
  orx   g00748(.a(n800), .b(n793), .O(n801));
  invx  g00749(.a(n801), .O(n802));
  andx  g00750(.a(n802), .b(n792), .O(n803));
  orx   g00751(.a(n803), .b(n68), .O(n804));
  andx  g00752(.a(n99), .b(pi10), .O(n805));
  invx  g00753(.a(n805), .O(n806));
  andx  g00754(.a(n806), .b(n804), .O(n807));
  andx  g00755(.a(n807), .b(n785), .O(n808));
  andx  g00756(.a(n808), .b(n783), .O(n809));
  andx  g00757(.a(n809), .b(n781), .O(n810));
  orx   g00758(.a(n330), .b(n47), .O(n811));
  andx  g00759(.a(n291), .b(pi06), .O(n812));
  invx  g00760(.a(n812), .O(n813));
  andx  g00761(.a(n813), .b(n811), .O(n814));
  andx  g00762(.a(n814), .b(n810), .O(n815));
  andx  g00763(.a(n815), .b(n779), .O(n816));
  orx   g00764(.a(n816), .b(n75), .O(n817));
  orx   g00765(.a(n115), .b(n79), .O(n818));
  invx  g00766(.a(n257), .O(n819));
  orx   g00767(.a(n819), .b(n46), .O(n820));
  andx  g00768(.a(n79), .b(n45), .O(n821));
  orx   g00769(.a(n821), .b(n78), .O(n822));
  orx   g00770(.a(n822), .b(n84), .O(n823));
  andx  g00771(.a(n823), .b(n820), .O(n824));
  andx  g00772(.a(n824), .b(n818), .O(n825));
  andx  g00773(.a(n825), .b(n817), .O(n826));
  invx  g00774(.a(n826), .O(n827));
  andx  g00775(.a(n827), .b(n604), .O(n828));
  andx  g00776(.a(n826), .b(n610), .O(n829));
  orx   g00777(.a(n829), .b(n828), .O(n830));
  orx   g00778(.a(n830), .b(n404), .O(n831));
  orx   g00779(.a(n831), .b(n777), .O(n832));
  orx   g00780(.a(n611), .b(n179), .O(n833));
  orx   g00781(.a(n826), .b(n610), .O(n834));
  orx   g00782(.a(n827), .b(n604), .O(n835));
  andx  g00783(.a(n835), .b(n834), .O(n836));
  andx  g00784(.a(n836), .b(n403), .O(n837));
  orx   g00785(.a(n837), .b(n833), .O(n838));
  andx  g00786(.a(n838), .b(n832), .O(n839));
  andx  g00787(.a(n554), .b(n214), .O(n840));
  invx  g00788(.a(n840), .O(n841));
  orx   g00789(.a(n607), .b(n612), .O(n842));
  andx  g00790(.a(n842), .b(n841), .O(n843));
  andx  g00791(.a(n613), .b(n606), .O(n844));
  andx  g00792(.a(n844), .b(n840), .O(n845));
  orx   g00793(.a(n845), .b(n843), .O(n846));
  andx  g00794(.a(n846), .b(n839), .O(n847));
  andx  g00795(.a(n837), .b(n833), .O(n848));
  andx  g00796(.a(n831), .b(n777), .O(n849));
  orx   g00797(.a(n849), .b(n848), .O(n850));
  orx   g00798(.a(n844), .b(n840), .O(n851));
  orx   g00799(.a(n842), .b(n841), .O(n852));
  andx  g00800(.a(n852), .b(n851), .O(n853));
  andx  g00801(.a(n853), .b(n850), .O(n854));
  orx   g00802(.a(n854), .b(n847), .O(n855));
  andx  g00803(.a(n617), .b(n626), .O(n856));
  andx  g00804(.a(n616), .b(n626), .O(n857));
  andx  g00805(.a(n617), .b(n616), .O(n858));
  orx   g00806(.a(n858), .b(n857), .O(n859));
  orx   g00807(.a(n859), .b(n856), .O(n860));
  andx  g00808(.a(n860), .b(n252), .O(n861));
  orx   g00809(.a(n618), .b(n615), .O(n862));
  orx   g00810(.a(n620), .b(n615), .O(n863));
  invx  g00811(.a(n858), .O(n864));
  andx  g00812(.a(n864), .b(n863), .O(n865));
  andx  g00813(.a(n865), .b(n862), .O(n866));
  andx  g00814(.a(n488), .b(n252), .O(n867));
  invx  g00815(.a(n867), .O(n868));
  andx  g00816(.a(n868), .b(n866), .O(n869));
  orx   g00817(.a(n869), .b(n861), .O(n870));
  andx  g00818(.a(n870), .b(n855), .O(n871));
  orx   g00819(.a(n853), .b(n850), .O(n872));
  orx   g00820(.a(n846), .b(n839), .O(n873));
  andx  g00821(.a(n873), .b(n872), .O(n874));
  orx   g00822(.a(n866), .b(n248), .O(n875));
  orx   g00823(.a(n867), .b(n860), .O(n876));
  andx  g00824(.a(n876), .b(n875), .O(n877));
  andx  g00825(.a(n877), .b(n874), .O(n878));
  orx   g00826(.a(n878), .b(n871), .O(n879));
  orx   g00827(.a(n879), .b(n776), .O(n880));
  orx   g00828(.a(n877), .b(n874), .O(n881));
  orx   g00829(.a(n870), .b(n855), .O(n882));
  andx  g00830(.a(n882), .b(n881), .O(n883));
  orx   g00831(.a(n883), .b(n775), .O(n884));
  andx  g00832(.a(n884), .b(n880), .O(n885));
  andx  g00833(.a(n379), .b(n338), .O(n890));
  invx  g00834(.a(n890), .O(n891));
  andx  g00835(.a(n675), .b(n586), .O(n892));
  invx  g00836(.a(n892), .O(n893));
  andx  g00837(.a(n682), .b(n592), .O(n894));
  orx   g00838(.a(n894), .b(n381), .O(n895));
  andx  g00839(.a(n895), .b(n893), .O(n896));
  orx   g00840(.a(n896), .b(n891), .O(n897));
  orx   g00841(.a(n675), .b(n586), .O(n898));
  andx  g00842(.a(n898), .b(n380), .O(n899));
  orx   g00843(.a(n899), .b(n892), .O(n900));
  orx   g00844(.a(n900), .b(n890), .O(n901));
  andx  g00845(.a(n901), .b(n897), .O(n902));
  andx  g00846(.a(n902), .b(n928), .O(n903));
  andx  g00847(.a(n900), .b(n890), .O(n906));
  andx  g00848(.a(n896), .b(n891), .O(n907));
  orx   g00849(.a(n907), .b(n906), .O(n908));
  andx  g00850(.a(n908), .b(n936), .O(n909));
  orx   g00851(.a(n909), .b(n903), .O(n910));
  orx   g00852(.a(n910), .b(n752), .O(n911));
  andx  g00853(.a(n910), .b(n752), .O(n912));
  invx  g00854(.a(n912), .O(n913));
  andx  g00855(.a(n913), .b(n911), .O(n914));
  andx  g00856(.a(n379), .b(n299), .O(n915));
  invx  g00857(.a(n915), .O(n916));
  andx  g00858(.a(n883), .b(n775), .O(n917));
  andx  g00859(.a(n879), .b(n776), .O(n918));
  orx   g00860(.a(n918), .b(n917), .O(n919));
  orx   g00861(.a(n765), .b(n919), .O(n923));
  andx  g00862(.a(n757), .b(n759), .O(n924));
  andx  g00863(.a(n763), .b(n753), .O(n925));
  orx   g00864(.a(n925), .b(n924), .O(n926));
  orx   g00865(.a(n926), .b(n885), .O(n927));
  andx  g00866(.a(n927), .b(n923), .O(n928));
  orx   g00867(.a(n928), .b(n900), .O(n929));
  orx   g00868(.a(n928), .b(n890), .O(n930));
  andx  g00869(.a(n930), .b(n901), .O(n931));
  andx  g00870(.a(n931), .b(n929), .O(n932));
  orx   g00871(.a(n932), .b(n916), .O(n933));
  andx  g00872(.a(n926), .b(n885), .O(n934));
  andx  g00873(.a(n765), .b(n919), .O(n935));
  orx   g00874(.a(n935), .b(n934), .O(n936));
  andx  g00875(.a(n936), .b(n896), .O(n937));
  andx  g00876(.a(n936), .b(n891), .O(n938));
  orx   g00877(.a(n938), .b(n907), .O(n939));
  orx   g00878(.a(n939), .b(n937), .O(n940));
  orx   g00879(.a(n940), .b(n915), .O(n941));
  andx  g00880(.a(n941), .b(n933), .O(n942));
  andx  g00881(.a(n499), .b(n376), .O(n943));
  andx  g00882(.a(n917), .b(n943), .O(n947));
  invx  g00883(.a(n943), .O(n948));
  andx  g00884(.a(n880), .b(n948), .O(n954));
  orx   g00885(.a(n954), .b(n947), .O(n955));
  andx  g00886(.a(n488), .b(n438), .O(n956));
  invx  g00887(.a(n956), .O(n957));
  andx  g00888(.a(n876), .b(n874), .O(n958));
  orx   g00889(.a(n958), .b(n861), .O(n959));
  andx  g00890(.a(n959), .b(n957), .O(n960));
  orx   g00891(.a(n869), .b(n855), .O(n961));
  andx  g00892(.a(n961), .b(n875), .O(n962));
  andx  g00893(.a(n962), .b(n956), .O(n963));
  orx   g00894(.a(n963), .b(n960), .O(n964));
  andx  g00895(.a(n835), .b(n403), .O(n969));
  invx  g00896(.a(n969), .O(n970));
  andx  g00897(.a(n836), .b(n250), .O(n971));
  andx  g00898(.a(n971), .b(n970), .O(n972));
  invx  g00899(.a(n971), .O(n973));
  andx  g00900(.a(n973), .b(n969), .O(n974));
  orx   g00901(.a(n974), .b(n972), .O(n975));
  andx  g00902(.a(n837), .b(n777), .O(n976));
  andx  g00903(.a(n605), .b(n214), .O(n977));
  andx  g00904(.a(n977), .b(n976), .O(n978));
  invx  g00905(.a(n978), .O(n979));
  orx   g00906(.a(n977), .b(n976), .O(n980));
  andx  g00907(.a(n980), .b(n979), .O(n981));
  orx   g00908(.a(n981), .b(n975), .O(n982));
  invx  g00909(.a(n975), .O(n983));
  invx  g00910(.a(n980), .O(n984));
  orx   g00911(.a(n984), .b(n978), .O(n985));
  orx   g00912(.a(n985), .b(n983), .O(n986));
  andx  g00913(.a(n986), .b(n982), .O(n987));
  orx   g00914(.a(n842), .b(n839), .O(n988));
  orx   g00915(.a(n841), .b(n839), .O(n989));
  andx  g00916(.a(n989), .b(n852), .O(n990));
  andx  g00917(.a(n990), .b(n988), .O(n991));
  orx   g00918(.a(n991), .b(n248), .O(n992));
  andx  g00919(.a(n844), .b(n850), .O(n993));
  andx  g00920(.a(n840), .b(n850), .O(n994));
  orx   g00921(.a(n994), .b(n845), .O(n995));
  orx   g00922(.a(n995), .b(n993), .O(n996));
  andx  g00923(.a(n554), .b(n252), .O(n997));
  orx   g00924(.a(n997), .b(n996), .O(n998));
  andx  g00925(.a(n998), .b(n992), .O(n999));
  orx   g00926(.a(n999), .b(n987), .O(n1000));
  andx  g00927(.a(n985), .b(n983), .O(n1001));
  orx   g00928(.a(n1150), .b(n1001), .O(n1003));
  andx  g00929(.a(n996), .b(n252), .O(n1004));
  invx  g00930(.a(n997), .O(n1005));
  andx  g00931(.a(n1005), .b(n991), .O(n1006));
  orx   g00932(.a(n1006), .b(n1004), .O(n1007));
  orx   g00933(.a(n1007), .b(n1003), .O(n1008));
  andx  g00934(.a(n1008), .b(n1000), .O(n1009));
  andx  g00935(.a(n1009), .b(n964), .O(n1010));
  orx   g00936(.a(n962), .b(n956), .O(n1011));
  orx   g00937(.a(n959), .b(n957), .O(n1012));
  andx  g00938(.a(n1012), .b(n1011), .O(n1013));
  andx  g00939(.a(n1007), .b(n1003), .O(n1014));
  andx  g00940(.a(n999), .b(n987), .O(n1015));
  orx   g00941(.a(n1015), .b(n1014), .O(n1016));
  andx  g00942(.a(n1016), .b(n1013), .O(n1017));
  orx   g00943(.a(n1017), .b(n1010), .O(n1018));
  orx   g00944(.a(n1018), .b(n955), .O(n1019));
  andx  g00945(.a(n1018), .b(n955), .O(n1020));
  invx  g00946(.a(n1020), .O(n1021));
  andx  g00947(.a(n1021), .b(n1019), .O(n1022));
  andx  g00948(.a(n885), .b(n757), .O(n1023));
  invx  g00949(.a(n1023), .O(n1024));
  andx  g00950(.a(n919), .b(n763), .O(n1025));
  orx   g00951(.a(n1025), .b(n759), .O(n1026));
  andx  g00952(.a(n1026), .b(n1024), .O(n1027));
  andx  g00953(.a(n338), .b(n255), .O(n1028));
  andx  g00954(.a(n1028), .b(n1027), .O(n1029));
  orx   g00955(.a(n885), .b(n757), .O(n1030));
  andx  g00956(.a(n1030), .b(n753), .O(n1031));
  orx   g00957(.a(n1031), .b(n1023), .O(n1032));
  invx  g00958(.a(n1028), .O(n1033));
  andx  g00959(.a(n1033), .b(n1032), .O(n1034));
  orx   g00960(.a(n1034), .b(n1029), .O(n1035));
  andx  g00961(.a(n1035), .b(n1022), .O(n1036));
  invx  g00962(.a(n1019), .O(n1037));
  orx   g00963(.a(n1020), .b(n1037), .O(n1038));
  orx   g00964(.a(n1033), .b(n1032), .O(n1039));
  orx   g00965(.a(n1028), .b(n1027), .O(n1040));
  andx  g00966(.a(n1040), .b(n1039), .O(n1041));
  andx  g00967(.a(n1041), .b(n1038), .O(n1042));
  orx   g00968(.a(n1042), .b(n1036), .O(n1043));
  orx   g00969(.a(n1043), .b(n942), .O(n1044));
  andx  g00970(.a(n940), .b(n915), .O(n1045));
  andx  g00971(.a(n932), .b(n916), .O(n1046));
  orx   g00972(.a(n1046), .b(n1045), .O(n1047));
  orx   g00973(.a(n1041), .b(n1038), .O(n1048));
  orx   g00974(.a(n1035), .b(n1022), .O(n1049));
  andx  g00975(.a(n1049), .b(n1048), .O(n1050));
  orx   g00976(.a(n1050), .b(n1047), .O(n1051));
  andx  g00977(.a(n1051), .b(n1044), .O(n1052));
  orx   g00978(.a(n908), .b(n936), .O(n1053));
  orx   g00979(.a(n902), .b(n928), .O(n1054));
  andx  g00980(.a(n1054), .b(n1053), .O(n1055));
  andx  g00981(.a(n1055), .b(n731), .O(n1056));
  invx  g00982(.a(n1056), .O(n1057));
  andx  g00983(.a(n910), .b(n750), .O(n1058));
  orx   g00984(.a(n1058), .b(n733), .O(n1059));
  andx  g00985(.a(n1059), .b(n1057), .O(n1060));
  andx  g00986(.a(n827), .b(n250), .O(n1061));
  invx  g00987(.a(n1061), .O(n1062));
  andx  g00988(.a(n1062), .b(n1060), .O(n1063));
  orx   g00989(.a(n1055), .b(n731), .O(n1064));
  andx  g00990(.a(n1064), .b(n300), .O(n1065));
  orx   g00991(.a(n1065), .b(n1056), .O(n1066));
  andx  g00992(.a(n1061), .b(n1066), .O(n1067));
  orx   g00993(.a(n1067), .b(n1063), .O(n1068));
  orx   g00994(.a(n1068), .b(n1052), .O(n1069));
  andx  g00995(.a(n1050), .b(n1047), .O(n1070));
  andx  g00996(.a(n1043), .b(n942), .O(n1071));
  orx   g00997(.a(n1071), .b(n1070), .O(n1072));
  orx   g00998(.a(n1061), .b(n1066), .O(n1073));
  orx   g00999(.a(n1062), .b(n1060), .O(n1074));
  andx  g01000(.a(n1074), .b(n1073), .O(n1075));
  orx   g01001(.a(n1075), .b(n1072), .O(n1076));
  andx  g01002(.a(n1076), .b(n1069), .O(n1077));
  andx  g01003(.a(n1077), .b(n914), .O(n1078));
  invx  g01004(.a(n914), .O(n1079));
  andx  g01005(.a(n1075), .b(n1072), .O(n1080));
  andx  g01006(.a(n1068), .b(n1052), .O(n1081));
  orx   g01007(.a(n1081), .b(n1080), .O(n1082));
  andx  g01008(.a(n1082), .b(n1079), .O(n1083));
  orx   g01009(.a(n1083), .b(n1078), .O(n1084));
  andx  g01010(.a(n1084), .b(n379), .O(n1085));
  andx  g01011(.a(n1085), .b(n914), .O(n1086));
  andx  g01012(.a(n1077), .b(n1079), .O(n1088));
  orx   g01013(.a(n1060), .b(n1072), .O(n1089));
  andx  g01014(.a(n1060), .b(n1072), .O(n1090));
  orx   g01015(.a(n1090), .b(n826), .O(n1091));
  andx  g01016(.a(n1091), .b(n1089), .O(n1092));
  andx  g01017(.a(n1092), .b(n250), .O(n1093));
  andx  g01018(.a(n827), .b(n379), .O(n1094));
  andx  g01019(.a(n932), .b(n915), .O(n1095));
  orx   g01020(.a(n932), .b(n915), .O(n1096));
  andx  g01021(.a(n1096), .b(n1050), .O(n1097));
  orx   g01022(.a(n1097), .b(n1095), .O(n1098));
  orx   g01023(.a(n1098), .b(n1094), .O(n1099));
  invx  g01024(.a(n1095), .O(n1100));
  andx  g01025(.a(n940), .b(n916), .O(n1101));
  orx   g01026(.a(n1101), .b(n1043), .O(n1102));
  andx  g01027(.a(n1102), .b(n1100), .O(n1103));
  orx   g01028(.a(n1103), .b(n826), .O(n1104));
  andx  g01029(.a(n1104), .b(n1099), .O(n1105));
  andx  g01030(.a(n299), .b(n255), .O(n1106));
  invx  g01031(.a(n1106), .O(n1107));
  andx  g01032(.a(n1033), .b(n1027), .O(n1108));
  andx  g01033(.a(n1028), .b(n1032), .O(n1109));
  invx  g01034(.a(n1109), .O(n1110));
  andx  g01035(.a(n1110), .b(n1038), .O(n1111));
  orx   g01036(.a(n1111), .b(n1108), .O(n1112));
  orx   g01037(.a(n1112), .b(n1107), .O(n1113));
  invx  g01038(.a(n1108), .O(n1114));
  orx   g01039(.a(n1109), .b(n1022), .O(n1115));
  andx  g01040(.a(n1115), .b(n1114), .O(n1116));
  orx   g01041(.a(n1116), .b(n1106), .O(n1117));
  andx  g01042(.a(n1117), .b(n1113), .O(n1118));
  andx  g01043(.a(n488), .b(n376), .O(n1119));
  invx  g01044(.a(n1119), .O(n1120));
  andx  g01045(.a(n959), .b(n956), .O(n1121));
  invx  g01046(.a(n1121), .O(n1122));
  andx  g01047(.a(n962), .b(n957), .O(n1123));
  orx   g01048(.a(n1123), .b(n1016), .O(n1124));
  andx  g01049(.a(n1124), .b(n1122), .O(n1125));
  andx  g01050(.a(n1125), .b(n1120), .O(n1126));
  invx  g01051(.a(n1126), .O(n1127));
  andx  g01052(.a(n554), .b(n438), .O(n1128));
  andx  g01053(.a(n998), .b(n987), .O(n1129));
  orx   g01054(.a(n1129), .b(n1004), .O(n1130));
  orx   g01055(.a(n1130), .b(n1128), .O(n1131));
  invx  g01056(.a(n1131), .O(n1132));
  andx  g01057(.a(n1130), .b(n1128), .O(n1133));
  orx   g01058(.a(n1133), .b(n1132), .O(n1134));
  andx  g01059(.a(n829), .b(n83), .O(n1135));
  andx  g01060(.a(n1135), .b(n403), .O(n1136));
  orx   g01061(.a(n1136), .b(n250), .O(n1137));
  invx  g01062(.a(n1137), .O(n1138));
  andx  g01063(.a(n836), .b(n214), .O(n1139));
  andx  g01064(.a(n971), .b(n403), .O(n1140));
  invx  g01065(.a(n1140), .O(n1141));
  andx  g01066(.a(n1141), .b(n1139), .O(n1142));
  invx  g01067(.a(n1139), .O(n1143));
  andx  g01068(.a(n1140), .b(n1143), .O(n1144));
  orx   g01069(.a(n1144), .b(n1142), .O(n1145));
  invx  g01070(.a(n1145), .O(n1146));
  andx  g01071(.a(n1146), .b(n1138), .O(n1147));
  andx  g01072(.a(n1145), .b(n1137), .O(n1148));
  orx   g01073(.a(n1148), .b(n1147), .O(n1149));
  andx  g01074(.a(n977), .b(n975), .O(n1150));
  orx   g01075(.a(n1150), .b(n978), .O(n1151));
  andx  g01076(.a(n1151), .b(n252), .O(n1152));
  andx  g01077(.a(n605), .b(n252), .O(n1153));
  orx   g01078(.a(n1153), .b(n1151), .O(n1154));
  invx  g01079(.a(n1154), .O(n1155));
  orx   g01080(.a(n1155), .b(n1152), .O(n1156));
  andx  g01081(.a(n1156), .b(n1149), .O(n1157));
  invx  g01082(.a(n1149), .O(n1158));
  invx  g01083(.a(n1152), .O(n1159));
  andx  g01084(.a(n1154), .b(n1159), .O(n1160));
  andx  g01085(.a(n1160), .b(n1158), .O(n1161));
  orx   g01086(.a(n1161), .b(n1157), .O(n1162));
  orx   g01087(.a(n1162), .b(n1134), .O(n1163));
  invx  g01088(.a(n1133), .O(n1164));
  andx  g01089(.a(n1164), .b(n1131), .O(n1165));
  orx   g01090(.a(n1160), .b(n1158), .O(n1166));
  orx   g01091(.a(n1156), .b(n1149), .O(n1167));
  andx  g01092(.a(n1167), .b(n1166), .O(n1168));
  orx   g01093(.a(n1168), .b(n1165), .O(n1169));
  andx  g01094(.a(n1169), .b(n1163), .O(n1170));
  andx  g01095(.a(n1170), .b(n1127), .O(n1171));
  andx  g01096(.a(n1168), .b(n1165), .O(n1172));
  andx  g01097(.a(n1162), .b(n1134), .O(n1173));
  orx   g01098(.a(n1173), .b(n1172), .O(n1174));
  andx  g01099(.a(n1174), .b(n1126), .O(n1175));
  orx   g01100(.a(n1175), .b(n1171), .O(n1176));
  orx   g01101(.a(n1016), .b(n1013), .O(n1177));
  orx   g01102(.a(n1009), .b(n964), .O(n1178));
  andx  g01103(.a(n1178), .b(n1177), .O(n1179));
  andx  g01104(.a(n1179), .b(n917), .O(n1180));
  orx   g01105(.a(n1179), .b(n917), .O(n1181));
  andx  g01106(.a(n1181), .b(n943), .O(n1182));
  orx   g01107(.a(n1182), .b(n1180), .O(n1183));
  andx  g01108(.a(n1183), .b(n338), .O(n1184));
  orx   g01109(.a(n1018), .b(n880), .O(n1185));
  andx  g01110(.a(n1018), .b(n880), .O(n1186));
  orx   g01111(.a(n1186), .b(n948), .O(n1187));
  andx  g01112(.a(n1187), .b(n1185), .O(n1188));
  andx  g01113(.a(n499), .b(n338), .O(n1189));
  invx  g01114(.a(n1189), .O(n1190));
  andx  g01115(.a(n1190), .b(n1188), .O(n1191));
  orx   g01116(.a(n1191), .b(n1184), .O(n1192));
  andx  g01117(.a(n1192), .b(n1176), .O(n1193));
  orx   g01118(.a(n1174), .b(n1126), .O(n1194));
  orx   g01119(.a(n1170), .b(n1127), .O(n1195));
  andx  g01120(.a(n1195), .b(n1194), .O(n1196));
  orx   g01121(.a(n1188), .b(n551), .O(n1197));
  orx   g01122(.a(n1189), .b(n1183), .O(n1198));
  andx  g01123(.a(n1198), .b(n1197), .O(n1199));
  andx  g01124(.a(n1199), .b(n1196), .O(n1200));
  orx   g01125(.a(n1200), .b(n1193), .O(n1201));
  orx   g01126(.a(n1201), .b(n1118), .O(n1202));
  andx  g01127(.a(n1116), .b(n1106), .O(n1203));
  andx  g01128(.a(n1112), .b(n1107), .O(n1204));
  orx   g01129(.a(n1204), .b(n1203), .O(n1205));
  orx   g01130(.a(n1199), .b(n1196), .O(n1206));
  orx   g01131(.a(n1192), .b(n1176), .O(n1207));
  andx  g01132(.a(n1207), .b(n1206), .O(n1208));
  orx   g01133(.a(n1208), .b(n1205), .O(n1209));
  andx  g01134(.a(n1209), .b(n1202), .O(n1210));
  orx   g01135(.a(n1210), .b(n1105), .O(n1211));
  invx  g01136(.a(n1094), .O(n1212));
  andx  g01137(.a(n1103), .b(n1212), .O(n1213));
  andx  g01138(.a(n1098), .b(n827), .O(n1214));
  orx   g01139(.a(n1214), .b(n1213), .O(n1215));
  andx  g01140(.a(n1208), .b(n1205), .O(n1216));
  andx  g01141(.a(n1201), .b(n1118), .O(n1217));
  orx   g01142(.a(n1217), .b(n1216), .O(n1218));
  orx   g01143(.a(n1218), .b(n1215), .O(n1219));
  andx  g01144(.a(n1219), .b(n1211), .O(n1220));
  andx  g01145(.a(n1220), .b(n1093), .O(n1221));
  andx  g01146(.a(n1066), .b(n1052), .O(n1222));
  orx   g01147(.a(n1066), .b(n1052), .O(n1223));
  andx  g01148(.a(n1223), .b(n827), .O(n1224));
  orx   g01149(.a(n1224), .b(n1222), .O(n1225));
  orx   g01150(.a(n1225), .b(n179), .O(n1226));
  andx  g01151(.a(n1218), .b(n1215), .O(n1227));
  andx  g01152(.a(n1210), .b(n1105), .O(n1228));
  orx   g01153(.a(n1228), .b(n1227), .O(n1229));
  andx  g01154(.a(n1229), .b(n1226), .O(n1230));
  orx   g01155(.a(n1230), .b(n1221), .O(n1231));
  andx  g01156(.a(n1231), .b(n1088), .O(n1232));
  invx  g01157(.a(n1088), .O(n1233));
  orx   g01158(.a(n1229), .b(n1226), .O(n1234));
  orx   g01159(.a(n1220), .b(n1093), .O(n1235));
  andx  g01160(.a(n1235), .b(n1234), .O(n1236));
  andx  g01161(.a(n1236), .b(n1233), .O(n1237));
  orx   g01162(.a(n1237), .b(n1232), .O(n1238));
  andx  g01163(.a(n1238), .b(n1580), .O(n1239));
  invx  g01164(.a(n1239), .O(n1240));
  andx  g01165(.a(n914), .b(n499), .O(n1241));
  invx  g01166(.a(n1241), .O(n1242));
  andx  g01167(.a(n1084), .b(n255), .O(n1243));
  invx  g01168(.a(n1243), .O(n1244));
  andx  g01169(.a(n1244), .b(n1242), .O(n1245));
  andx  g01170(.a(n1243), .b(n1241), .O(n1246));
  orx   g01171(.a(n1246), .b(n1245), .O(n1247));
  invx  g01172(.a(n1580), .O(n1248));
  orx   g01173(.a(n1236), .b(n1233), .O(n1249));
  orx   g01174(.a(n1231), .b(n1088), .O(n1250));
  andx  g01175(.a(n1250), .b(n1249), .O(n1251));
  orx   g01176(.a(n1251), .b(n378), .O(n1252));
  andx  g01177(.a(n1252), .b(n1248), .O(n1253));
  orx   g01178(.a(n1253), .b(n1247), .O(n1254));
  andx  g01179(.a(n1254), .b(n1240), .O(n1255));
  andx  g01180(.a(n1236), .b(n1088), .O(n1256));
  invx  g01181(.a(n1256), .O(n1257));
  andx  g01182(.a(n1220), .b(n1092), .O(n1258));
  orx   g01183(.a(n1258), .b(n179), .O(n1259));
  andx  g01184(.a(n1218), .b(n1099), .O(n1260));
  orx   g01185(.a(n1260), .b(n1214), .O(n1261));
  orx   g01186(.a(n1261), .b(n378), .O(n1262));
  andx  g01187(.a(n488), .b(n338), .O(n1263));
  invx  g01188(.a(n1263), .O(n1264));
  orx   g01189(.a(n1171), .b(n1264), .O(n1267));
  orx   g01190(.a(n1194), .b(n1263), .O(n1269));
  andx  g01191(.a(n1269), .b(n1267), .O(n1270));
  andx  g01192(.a(n605), .b(n438), .O(n1271));
  invx  g01193(.a(n1271), .O(n1272));
  orx   g01194(.a(n1155), .b(n1149), .O(n1273));
  andx  g01195(.a(n1273), .b(n1159), .O(n1274));
  andx  g01196(.a(n1274), .b(n1272), .O(n1275));
  orx   g01197(.a(n1274), .b(n1272), .O(n1276));
  invx  g01198(.a(n1276), .O(n1277));
  orx   g01199(.a(n1277), .b(n1275), .O(n1278));
  andx  g01200(.a(n1141), .b(n1143), .O(n1279));
  orx   g01201(.a(n1279), .b(n1138), .O(n1280));
  invx  g01202(.a(n1280), .O(n1281));
  andx  g01203(.a(n1281), .b(n252), .O(n1282));
  invx  g01204(.a(n1282), .O(n1283));
  andx  g01205(.a(n836), .b(n252), .O(n1284));
  orx   g01206(.a(n1284), .b(n1281), .O(n1285));
  andx  g01207(.a(n1285), .b(n1283), .O(n1286));
  invx  g01208(.a(n1286), .O(n1287));
  andx  g01209(.a(n1287), .b(n214), .O(n1288));
  andx  g01210(.a(n1286), .b(n215), .O(n1289));
  orx   g01211(.a(n1289), .b(n1288), .O(n1290));
  invx  g01212(.a(n1290), .O(n1291));
  orx   g01213(.a(n1291), .b(n1278), .O(n1292));
  invx  g01214(.a(n1275), .O(n1293));
  andx  g01215(.a(n1276), .b(n1293), .O(n1294));
  orx   g01216(.a(n1290), .b(n1294), .O(n1295));
  andx  g01217(.a(n1295), .b(n1292), .O(n1296));
  andx  g01218(.a(n554), .b(n376), .O(n1297));
  orx   g01219(.a(n1162), .b(n1132), .O(n1298));
  andx  g01220(.a(n1298), .b(n1164), .O(n1299));
  orx   g01221(.a(n1299), .b(n1297), .O(n1300));
  invx  g01222(.a(n1297), .O(n1301));
  andx  g01223(.a(n1168), .b(n1131), .O(n1302));
  orx   g01224(.a(n1302), .b(n1133), .O(n1303));
  orx   g01225(.a(n1303), .b(n1301), .O(n1304));
  andx  g01226(.a(n1304), .b(n1300), .O(n1305));
  orx   g01227(.a(n1305), .b(n1296), .O(n1306));
  andx  g01228(.a(n1290), .b(n1294), .O(n1307));
  andx  g01229(.a(n1291), .b(n1278), .O(n1308));
  orx   g01230(.a(n1308), .b(n1307), .O(n1309));
  andx  g01231(.a(n1303), .b(n1301), .O(n1310));
  andx  g01232(.a(n1299), .b(n1297), .O(n1311));
  orx   g01233(.a(n1311), .b(n1310), .O(n1312));
  orx   g01234(.a(n1312), .b(n1309), .O(n1313));
  andx  g01235(.a(n1313), .b(n1306), .O(n1314));
  andx  g01236(.a(n1314), .b(n1270), .O(n1315));
  andx  g01237(.a(n1194), .b(n1263), .O(n1316));
  andx  g01238(.a(n1171), .b(n1264), .O(n1317));
  orx   g01239(.a(n1317), .b(n1316), .O(n1318));
  andx  g01240(.a(n1312), .b(n1309), .O(n1319));
  andx  g01241(.a(n1305), .b(n1296), .O(n1320));
  orx   g01242(.a(n1320), .b(n1319), .O(n1321));
  andx  g01243(.a(n1321), .b(n1318), .O(n1322));
  orx   g01244(.a(n1322), .b(n1315), .O(n1323));
  andx  g01245(.a(n499), .b(n299), .O(n1324));
  invx  g01246(.a(n1324), .O(n1325));
  andx  g01247(.a(n1198), .b(n1196), .O(n1326));
  orx   g01248(.a(n1326), .b(n1184), .O(n1327));
  andx  g01249(.a(n1327), .b(n1325), .O(n1328));
  orx   g01250(.a(n1327), .b(n1325), .O(n1329));
  invx  g01251(.a(n1329), .O(n1330));
  orx   g01252(.a(n1330), .b(n1328), .O(n1331));
  andx  g01253(.a(n1331), .b(n1323), .O(n1332));
  orx   g01254(.a(n1321), .b(n1318), .O(n1333));
  orx   g01255(.a(n1314), .b(n1270), .O(n1334));
  andx  g01256(.a(n1334), .b(n1333), .O(n1335));
  invx  g01257(.a(n1328), .O(n1336));
  andx  g01258(.a(n1329), .b(n1336), .O(n1337));
  andx  g01259(.a(n1337), .b(n1335), .O(n1338));
  orx   g01260(.a(n1338), .b(n1332), .O(n1339));
  andx  g01261(.a(n827), .b(n255), .O(n1340));
  invx  g01262(.a(n1340), .O(n1341));
  andx  g01263(.a(n1208), .b(n1116), .O(n1342));
  orx   g01264(.a(n1208), .b(n1116), .O(n1343));
  andx  g01265(.a(n1343), .b(n1106), .O(n1344));
  orx   g01266(.a(n1344), .b(n1342), .O(n1345));
  andx  g01267(.a(n1345), .b(n1341), .O(n1346));
  orx   g01268(.a(n1201), .b(n1112), .O(n1347));
  andx  g01269(.a(n1201), .b(n1112), .O(n1348));
  orx   g01270(.a(n1348), .b(n1107), .O(n1349));
  andx  g01271(.a(n1349), .b(n1347), .O(n1350));
  andx  g01272(.a(n1350), .b(n1340), .O(n1351));
  orx   g01273(.a(n1351), .b(n1346), .O(n1352));
  andx  g01274(.a(n1352), .b(n1339), .O(n1353));
  orx   g01275(.a(n1337), .b(n1335), .O(n1354));
  orx   g01276(.a(n1331), .b(n1323), .O(n1355));
  andx  g01277(.a(n1355), .b(n1354), .O(n1356));
  orx   g01278(.a(n1350), .b(n1340), .O(n1357));
  orx   g01279(.a(n1345), .b(n1341), .O(n1358));
  andx  g01280(.a(n1358), .b(n1357), .O(n1359));
  andx  g01281(.a(n1359), .b(n1356), .O(n1360));
  orx   g01282(.a(n1360), .b(n1353), .O(n1361));
  orx   g01283(.a(n1361), .b(n1262), .O(n1362));
  orx   g01284(.a(n1210), .b(n1213), .O(n1363));
  andx  g01285(.a(n1363), .b(n1104), .O(n1364));
  andx  g01286(.a(n1364), .b(n379), .O(n1365));
  orx   g01287(.a(n1359), .b(n1356), .O(n1366));
  orx   g01288(.a(n1352), .b(n1339), .O(n1367));
  andx  g01289(.a(n1367), .b(n1366), .O(n1368));
  orx   g01290(.a(n1368), .b(n1365), .O(n1369));
  andx  g01291(.a(n1369), .b(n1362), .O(n1370));
  orx   g01292(.a(n1370), .b(n1259), .O(n1371));
  invx  g01293(.a(n1259), .O(n1372));
  andx  g01294(.a(n1368), .b(n1365), .O(n1373));
  andx  g01295(.a(n1361), .b(n1262), .O(n1374));
  orx   g01296(.a(n1374), .b(n1373), .O(n1375));
  orx   g01297(.a(n1375), .b(n1372), .O(n1376));
  andx  g01298(.a(n1376), .b(n1371), .O(n1377));
  andx  g01299(.a(n1377), .b(n1257), .O(n1378));
  andx  g01300(.a(n1375), .b(n1372), .O(n1379));
  andx  g01301(.a(n1370), .b(n1259), .O(n1380));
  orx   g01302(.a(n1380), .b(n1379), .O(n1381));
  andx  g01303(.a(n1381), .b(n1256), .O(n1382));
  orx   g01304(.a(n1382), .b(n1378), .O(n1383));
  andx  g01305(.a(n1383), .b(n379), .O(n1384));
  andx  g01306(.a(n1384), .b(n1255), .O(n1385));
  invx  g01307(.a(n1247), .O(n1386));
  andx  g01308(.a(n1238), .b(n379), .O(n1387));
  orx   g01309(.a(n1387), .b(n1580), .O(n1388));
  andx  g01310(.a(n1388), .b(n1386), .O(n1389));
  orx   g01311(.a(n1389), .b(n1239), .O(n1390));
  orx   g01312(.a(n1381), .b(n1256), .O(n1391));
  orx   g01313(.a(n1377), .b(n1257), .O(n1392));
  andx  g01314(.a(n1392), .b(n1391), .O(n1393));
  orx   g01315(.a(n1393), .b(n378), .O(n1394));
  andx  g01316(.a(n1394), .b(n1390), .O(n1395));
  orx   g01317(.a(n1395), .b(n1385), .O(n1396));
  invx  g01318(.a(n1246), .O(n1397));
  andx  g01319(.a(n1238), .b(n255), .O(n1398));
  andx  g01320(.a(n1398), .b(n1397), .O(n1399));
  orx   g01321(.a(n1251), .b(n254), .O(n1400));
  andx  g01322(.a(n1400), .b(n1246), .O(n1401));
  orx   g01323(.a(n1401), .b(n1399), .O(n1402));
  andx  g01324(.a(n914), .b(n488), .O(n1403));
  invx  g01325(.a(n1403), .O(n1404));
  orx   g01326(.a(n1082), .b(n1079), .O(n1405));
  orx   g01327(.a(n1077), .b(n914), .O(n1406));
  andx  g01328(.a(n1406), .b(n1405), .O(n1407));
  orx   g01329(.a(n1407), .b(n481), .O(n1408));
  andx  g01330(.a(n1408), .b(n1404), .O(n1409));
  andx  g01331(.a(n1084), .b(n499), .O(n1410));
  andx  g01332(.a(n1410), .b(n1403), .O(n1411));
  orx   g01333(.a(n1411), .b(n1409), .O(n1412));
  orx   g01334(.a(n1730), .b(n1402), .O(n1414));
  orx   g01335(.a(n1400), .b(n1246), .O(n1415));
  orx   g01336(.a(n1398), .b(n1397), .O(n1416));
  andx  g01337(.a(n1416), .b(n1415), .O(n1417));
  orx   g01338(.a(n1412), .b(n1417), .O(n1418));
  andx  g01339(.a(n1418), .b(n1414), .O(n1419));
  andx  g01340(.a(n1419), .b(n1396), .O(n1420));
  orx   g01341(.a(n1394), .b(n1390), .O(n1421));
  orx   g01342(.a(n1384), .b(n1255), .O(n1422));
  andx  g01343(.a(n1422), .b(n1421), .O(n1423));
  andx  g01344(.a(n1412), .b(n1417), .O(n1424));
  andx  g01345(.a(n1730), .b(n1402), .O(n1425));
  orx   g01346(.a(n1425), .b(n1424), .O(n1426));
  andx  g01347(.a(n1426), .b(n1423), .O(n1427));
  orx   g01348(.a(n1427), .b(n1420), .O(n1428));
  andx  g01349(.a(n1377), .b(n1256), .O(n1429));
  orx   g01350(.a(n1361), .b(n378), .O(n1430));
  andx  g01351(.a(n1430), .b(n1364), .O(n1431));
  andx  g01352(.a(n488), .b(n299), .O(n1432));
  invx  g01353(.a(n1432), .O(n1433));
  andx  g01354(.a(n1321), .b(n1263), .O(n1434));
  invx  g01355(.a(n1434), .O(n1435));
  andx  g01356(.a(n1314), .b(n1264), .O(n1436));
  orx   g01357(.a(n1436), .b(n1194), .O(n1437));
  andx  g01358(.a(n1437), .b(n1435), .O(n1438));
  orx   g01359(.a(n1438), .b(n1433), .O(n1439));
  orx   g01360(.a(n1321), .b(n1263), .O(n1440));
  andx  g01361(.a(n1440), .b(n1171), .O(n1441));
  orx   g01362(.a(n1441), .b(n1434), .O(n1442));
  orx   g01363(.a(n1442), .b(n1432), .O(n1443));
  andx  g01364(.a(n1443), .b(n1439), .O(n1444));
  andx  g01365(.a(n476), .b(n338), .O(n1445));
  invx  g01366(.a(n1445), .O(n1446));
  andx  g01367(.a(n1303), .b(n1296), .O(n1447));
  invx  g01368(.a(n1447), .O(n1448));
  andx  g01369(.a(n1299), .b(n1309), .O(n1449));
  orx   g01370(.a(n1449), .b(n1301), .O(n1450));
  andx  g01371(.a(n1450), .b(n1448), .O(n1451));
  andx  g01372(.a(n1451), .b(n1446), .O(n1452));
  andx  g01373(.a(n1285), .b(n214), .O(n1453));
  orx   g01374(.a(n1453), .b(n1282), .O(n1454));
  invx  g01375(.a(n1454), .O(n1455));
  andx  g01376(.a(n836), .b(n438), .O(n1456));
  andx  g01377(.a(n1456), .b(n248), .O(n1457));
  invx  g01378(.a(n1456), .O(n1458));
  andx  g01379(.a(n1458), .b(n252), .O(n1459));
  orx   g01380(.a(n1459), .b(n1457), .O(n1460));
  andx  g01381(.a(n1460), .b(n1455), .O(n1461));
  invx  g01382(.a(n1461), .O(n1462));
  orx   g01383(.a(n1460), .b(n1455), .O(n1463));
  andx  g01384(.a(n1463), .b(n1462), .O(n1464));
  invx  g01385(.a(n1464), .O(n1465));
  andx  g01386(.a(n605), .b(n376), .O(n1466));
  invx  g01387(.a(n1466), .O(n1467));
  andx  g01388(.a(n1290), .b(n1293), .O(n1468));
  orx   g01389(.a(n1468), .b(n1277), .O(n1469));
  andx  g01390(.a(n1469), .b(n1467), .O(n1470));
  invx  g01391(.a(n1470), .O(n1471));
  orx   g01392(.a(n1469), .b(n1467), .O(n1472));
  andx  g01393(.a(n1472), .b(n1471), .O(n1473));
  orx   g01394(.a(n1473), .b(n1465), .O(n1474));
  invx  g01395(.a(n1472), .O(n1475));
  orx   g01396(.a(n1475), .b(n1470), .O(n1476));
  orx   g01397(.a(n1476), .b(n1464), .O(n1477));
  andx  g01398(.a(n1477), .b(n1474), .O(n1478));
  orx   g01399(.a(n1478), .b(n1452), .O(n1479));
  orx   g01400(.a(n1303), .b(n1296), .O(n1480));
  andx  g01401(.a(n1480), .b(n1297), .O(n1481));
  orx   g01402(.a(n1481), .b(n1447), .O(n1482));
  orx   g01403(.a(n1482), .b(n1445), .O(n1483));
  andx  g01404(.a(n1476), .b(n1464), .O(n1484));
  andx  g01405(.a(n1473), .b(n1465), .O(n1485));
  orx   g01406(.a(n1485), .b(n1484), .O(n1486));
  orx   g01407(.a(n1486), .b(n1483), .O(n1487));
  andx  g01408(.a(n1487), .b(n1479), .O(n1488));
  andx  g01409(.a(n1488), .b(n1444), .O(n1489));
  andx  g01410(.a(n1442), .b(n1432), .O(n1490));
  andx  g01411(.a(n1438), .b(n1433), .O(n1491));
  orx   g01412(.a(n1491), .b(n1490), .O(n1492));
  andx  g01413(.a(n1486), .b(n1483), .O(n1493));
  andx  g01414(.a(n1478), .b(n1452), .O(n1494));
  orx   g01415(.a(n1494), .b(n1493), .O(n1495));
  andx  g01416(.a(n1495), .b(n1492), .O(n1496));
  orx   g01417(.a(n1496), .b(n1489), .O(n1497));
  andx  g01418(.a(n1327), .b(n1335), .O(n1498));
  orx   g01419(.a(n1327), .b(n1335), .O(n1499));
  andx  g01420(.a(n1499), .b(n1324), .O(n1500));
  orx   g01421(.a(n1500), .b(n1498), .O(n1501));
  andx  g01422(.a(n1501), .b(n827), .O(n1502));
  invx  g01423(.a(n1498), .O(n1503));
  invx  g01424(.a(n1327), .O(n1504));
  andx  g01425(.a(n1504), .b(n1323), .O(n1505));
  orx   g01426(.a(n1505), .b(n1325), .O(n1506));
  andx  g01427(.a(n1506), .b(n1503), .O(n1507));
  andx  g01428(.a(n827), .b(n499), .O(n1508));
  invx  g01429(.a(n1508), .O(n1509));
  andx  g01430(.a(n1509), .b(n1507), .O(n1510));
  orx   g01431(.a(n1510), .b(n1502), .O(n1511));
  andx  g01432(.a(n1511), .b(n1497), .O(n1512));
  orx   g01433(.a(n1495), .b(n1492), .O(n1513));
  orx   g01434(.a(n1488), .b(n1444), .O(n1514));
  andx  g01435(.a(n1514), .b(n1513), .O(n1515));
  orx   g01436(.a(n1507), .b(n826), .O(n1516));
  orx   g01437(.a(n1508), .b(n1501), .O(n1517));
  andx  g01438(.a(n1517), .b(n1516), .O(n1518));
  andx  g01439(.a(n1518), .b(n1515), .O(n1519));
  orx   g01440(.a(n1519), .b(n1512), .O(n1520));
  andx  g01441(.a(n1350), .b(n1341), .O(n1521));
  orx   g01442(.a(n1350), .b(n1341), .O(n1522));
  andx  g01443(.a(n1522), .b(n1356), .O(n1523));
  orx   g01444(.a(n1523), .b(n1521), .O(n1524));
  andx  g01445(.a(n1524), .b(n255), .O(n1525));
  orx   g01446(.a(n1525), .b(n1520), .O(n1526));
  orx   g01447(.a(n1518), .b(n1515), .O(n1527));
  orx   g01448(.a(n1511), .b(n1497), .O(n1528));
  andx  g01449(.a(n1528), .b(n1527), .O(n1529));
  invx  g01450(.a(n1521), .O(n1530));
  andx  g01451(.a(n1345), .b(n1340), .O(n1531));
  orx   g01452(.a(n1531), .b(n1339), .O(n1532));
  andx  g01453(.a(n1532), .b(n1530), .O(n1533));
  orx   g01454(.a(n1533), .b(n254), .O(n1534));
  orx   g01455(.a(n1534), .b(n1529), .O(n1535));
  andx  g01456(.a(n1535), .b(n1526), .O(n1536));
  orx   g01457(.a(n1536), .b(n1431), .O(n1537));
  andx  g01458(.a(n1368), .b(n379), .O(n1538));
  orx   g01459(.a(n1538), .b(n1261), .O(n1539));
  andx  g01460(.a(n1534), .b(n1529), .O(n1540));
  andx  g01461(.a(n1525), .b(n1520), .O(n1541));
  orx   g01462(.a(n1541), .b(n1540), .O(n1542));
  orx   g01463(.a(n1542), .b(n1539), .O(n1543));
  andx  g01464(.a(n1543), .b(n1537), .O(n1544));
  andx  g01465(.a(n1370), .b(n1372), .O(n1545));
  orx   g01466(.a(n1545), .b(n1544), .O(n1546));
  andx  g01467(.a(n1542), .b(n1539), .O(n1547));
  andx  g01468(.a(n1536), .b(n1431), .O(n1548));
  orx   g01469(.a(n1548), .b(n1547), .O(n1549));
  invx  g01470(.a(n1545), .O(n1550));
  orx   g01471(.a(n1550), .b(n1549), .O(n1551));
  andx  g01472(.a(n1551), .b(n1546), .O(n1552));
  andx  g01473(.a(n1552), .b(n1429), .O(n1553));
  invx  g01474(.a(n1429), .O(n1554));
  andx  g01475(.a(n1550), .b(n1549), .O(n1555));
  andx  g01476(.a(n1545), .b(n1544), .O(n1556));
  orx   g01477(.a(n1556), .b(n1555), .O(n1557));
  andx  g01478(.a(n1557), .b(n1554), .O(n1558));
  orx   g01479(.a(n1558), .b(n1553), .O(n1559));
  andx  g01480(.a(n1559), .b(n250), .O(n1560));
  invx  g01481(.a(n1560), .O(n1561));
  andx  g01482(.a(n1561), .b(n1428), .O(n1562));
  invx  g01483(.a(n1562), .O(n1563));
  orx   g01484(.a(n1426), .b(n1423), .O(n1564));
  orx   g01485(.a(n1419), .b(n1396), .O(n1565));
  andx  g01486(.a(n1565), .b(n1564), .O(n1566));
  andx  g01487(.a(n1560), .b(n1566), .O(n1567));
  andx  g01488(.a(n1388), .b(n1240), .O(n1568));
  orx   g01489(.a(n1568), .b(n1247), .O(n1569));
  invx  g01490(.a(n1569), .O(n1570));
  andx  g01491(.a(n1568), .b(n1247), .O(n1571));
  orx   g01492(.a(n1571), .b(n1570), .O(n1572));
  andx  g01493(.a(n1383), .b(n250), .O(n1573));
  andx  g01494(.a(n1573), .b(n1572), .O(n1574));
  orx   g01495(.a(n1572), .b(n1383), .O(n1575));
  invx  g01496(.a(n1085), .O(n1576));
  andx  g01497(.a(n914), .b(n255), .O(n1577));
  invx  g01498(.a(n1577), .O(n1578));
  andx  g01499(.a(n1578), .b(n1576), .O(n1579));
  andx  g01500(.a(n1577), .b(n1085), .O(n1580));
  orx   g01501(.a(n1580), .b(n1579), .O(n1581));
  invx  g01502(.a(n1581), .O(n1582));
  andx  g01503(.a(n1582), .b(n1086), .O(n1583));
  orx   g01504(.a(n1583), .b(n1238), .O(n1584));
  orx   g01505(.a(n1579), .b(n179), .O(n1587));
  invx  g01506(.a(n1587), .O(n1588));
  andx  g01507(.a(n1588), .b(n1584), .O(n1589));
  andx  g01508(.a(n1589), .b(n1575), .O(n1590));
  orx   g01509(.a(n1590), .b(n1574), .O(n1591));
  orx   g01510(.a(n1591), .b(n1567), .O(n1592));
  andx  g01511(.a(n1592), .b(n1563), .O(n1593));
  andx  g01512(.a(n1557), .b(n1429), .O(n1594));
  invx  g01513(.a(n1594), .O(n1595));
  andx  g01514(.a(n1517), .b(n1515), .O(n1596));
  orx   g01515(.a(n1596), .b(n1502), .O(n1597));
  orx   g01516(.a(n1597), .b(n481), .O(n1598));
  andx  g01517(.a(n554), .b(n299), .O(n1601));
  andx  g01518(.a(n1601), .b(n1479), .O(n1602));
  invx  g01519(.a(n1601), .O(n1603));
  andx  g01520(.a(n1603), .b(n1493), .O(n1604));
  orx   g01521(.a(n1604), .b(n1602), .O(n1605));
  invx  g01522(.a(n1605), .O(n1606));
  andx  g01523(.a(n1456), .b(n1454), .O(n1607));
  invx  g01524(.a(n1607), .O(n1608));
  andx  g01525(.a(n1458), .b(n1455), .O(n1609));
  orx   g01526(.a(n1609), .b(n248), .O(n1610));
  andx  g01527(.a(n1610), .b(n1608), .O(n1611));
  andx  g01528(.a(n1611), .b(n474), .O(n1612));
  invx  g01529(.a(n1612), .O(n1613));
  orx   g01530(.a(n1611), .b(n474), .O(n1614));
  andx  g01531(.a(n1614), .b(n1613), .O(n1615));
  andx  g01532(.a(n836), .b(n376), .O(n1616));
  invx  g01533(.a(n1616), .O(n1617));
  andx  g01534(.a(n1617), .b(n1615), .O(n1618));
  invx  g01535(.a(n1618), .O(n1619));
  orx   g01536(.a(n1617), .b(n1615), .O(n1620));
  andx  g01537(.a(n1620), .b(n1619), .O(n1621));
  invx  g01538(.a(n1621), .O(n1622));
  andx  g01539(.a(n338), .b(n602), .O(n1623));
  andx  g01540(.a(n1469), .b(n1465), .O(n1624));
  invx  g01541(.a(n1624), .O(n1625));
  invx  g01542(.a(n1469), .O(n1626));
  andx  g01543(.a(n1626), .b(n1464), .O(n1627));
  orx   g01544(.a(n1627), .b(n1467), .O(n1628));
  andx  g01545(.a(n1628), .b(n1625), .O(n1629));
  orx   g01546(.a(n1629), .b(n1623), .O(n1630));
  andx  g01547(.a(n1629), .b(n1623), .O(n1631));
  invx  g01548(.a(n1631), .O(n1632));
  andx  g01549(.a(n1632), .b(n1630), .O(n1633));
  orx   g01550(.a(n1633), .b(n1622), .O(n1634));
  invx  g01551(.a(n1634), .O(n1635));
  andx  g01552(.a(n1633), .b(n1622), .O(n1636));
  orx   g01553(.a(n1636), .b(n1635), .O(n1637));
  andx  g01554(.a(n1637), .b(n1606), .O(n1638));
  invx  g01555(.a(n1636), .O(n1639));
  andx  g01556(.a(n1639), .b(n1634), .O(n1640));
  andx  g01557(.a(n1640), .b(n1605), .O(n1641));
  orx   g01558(.a(n1641), .b(n1638), .O(n1642));
  andx  g01559(.a(n1488), .b(n1442), .O(n1643));
  invx  g01560(.a(n1643), .O(n1644));
  andx  g01561(.a(n1495), .b(n1438), .O(n1645));
  orx   g01562(.a(n1645), .b(n1433), .O(n1646));
  andx  g01563(.a(n1646), .b(n1644), .O(n1647));
  orx   g01564(.a(n1647), .b(n826), .O(n1648));
  orx   g01565(.a(n1488), .b(n1442), .O(n1649));
  andx  g01566(.a(n1649), .b(n1432), .O(n1650));
  orx   g01567(.a(n1650), .b(n1643), .O(n1651));
  andx  g01568(.a(n827), .b(n488), .O(n1652));
  orx   g01569(.a(n1652), .b(n1651), .O(n1653));
  andx  g01570(.a(n1653), .b(n1648), .O(n1654));
  orx   g01571(.a(n1654), .b(n1642), .O(n1655));
  orx   g01572(.a(n1640), .b(n1605), .O(n1656));
  orx   g01573(.a(n1637), .b(n1606), .O(n1657));
  andx  g01574(.a(n1657), .b(n1656), .O(n1658));
  andx  g01575(.a(n1651), .b(n827), .O(n1659));
  invx  g01576(.a(n1652), .O(n1660));
  andx  g01577(.a(n1660), .b(n1647), .O(n1661));
  orx   g01578(.a(n1661), .b(n1659), .O(n1662));
  orx   g01579(.a(n1662), .b(n1658), .O(n1663));
  andx  g01580(.a(n1663), .b(n1655), .O(n1664));
  andx  g01581(.a(n1664), .b(n1598), .O(n1665));
  invx  g01582(.a(n1598), .O(n1666));
  andx  g01583(.a(n1662), .b(n1658), .O(n1667));
  andx  g01584(.a(n1654), .b(n1642), .O(n1668));
  orx   g01585(.a(n1668), .b(n1667), .O(n1669));
  andx  g01586(.a(n1669), .b(n1666), .O(n1670));
  orx   g01587(.a(n1670), .b(n1665), .O(n1671));
  andx  g01588(.a(n1524), .b(n1520), .O(n1672));
  orx   g01589(.a(n1672), .b(n254), .O(n1673));
  invx  g01590(.a(n1673), .O(n1674));
  orx   g01591(.a(n1674), .b(n1671), .O(n1675));
  orx   g01592(.a(n1669), .b(n1666), .O(n1676));
  orx   g01593(.a(n1664), .b(n1598), .O(n1677));
  andx  g01594(.a(n1677), .b(n1676), .O(n1678));
  orx   g01595(.a(n1673), .b(n1678), .O(n1679));
  andx  g01596(.a(n1679), .b(n1675), .O(n1680));
  andx  g01597(.a(n1680), .b(n1547), .O(n1681));
  andx  g01598(.a(n1673), .b(n1678), .O(n1682));
  andx  g01599(.a(n1674), .b(n1671), .O(n1683));
  orx   g01600(.a(n1683), .b(n1682), .O(n1684));
  andx  g01601(.a(n1684), .b(n1537), .O(n1685));
  orx   g01602(.a(n1685), .b(n1681), .O(n1686));
  andx  g01603(.a(n1686), .b(n1551), .O(n1687));
  orx   g01604(.a(n1684), .b(n1537), .O(n1688));
  orx   g01605(.a(n1680), .b(n1547), .O(n1689));
  andx  g01606(.a(n1689), .b(n1688), .O(n1690));
  orx   g01607(.a(n1825), .b(n1687), .O(n1692));
  andx  g01608(.a(n1692), .b(n1595), .O(n1693));
  orx   g01609(.a(n1690), .b(n1556), .O(n1694));
  orx   g01610(.a(n1686), .b(n1551), .O(n1695));
  andx  g01611(.a(n1695), .b(n1694), .O(n1696));
  andx  g01612(.a(n1696), .b(n1594), .O(n1697));
  orx   g01613(.a(n1697), .b(n1693), .O(n1698));
  andx  g01614(.a(n1698), .b(n250), .O(n1699));
  andx  g01615(.a(n1699), .b(n1593), .O(n1700));
  orx   g01616(.a(n1561), .b(n1428), .O(n1701));
  invx  g01617(.a(n1574), .O(n1702));
  invx  g01618(.a(n1571), .O(n1703));
  andx  g01619(.a(n1703), .b(n1569), .O(n1704));
  andx  g01620(.a(n1704), .b(n1393), .O(n1705));
  invx  g01621(.a(n1589), .O(n1706));
  orx   g01622(.a(n1706), .b(n1705), .O(n1707));
  andx  g01623(.a(n1707), .b(n1702), .O(n1708));
  andx  g01624(.a(n1708), .b(n1701), .O(n1709));
  orx   g01625(.a(n1709), .b(n1562), .O(n1710));
  invx  g01626(.a(n1699), .O(n1711));
  andx  g01627(.a(n1711), .b(n1710), .O(n1712));
  orx   g01628(.a(n1712), .b(n1700), .O(n1713));
  andx  g01629(.a(n1559), .b(n379), .O(n1714));
  andx  g01630(.a(n1419), .b(n1390), .O(n1715));
  orx   g01631(.a(n1419), .b(n1390), .O(n1716));
  andx  g01632(.a(n1716), .b(n1384), .O(n1717));
  orx   g01633(.a(n1717), .b(n1715), .O(n1718));
  andx  g01634(.a(n1718), .b(n1714), .O(n1719));
  invx  g01635(.a(n1714), .O(n1720));
  orx   g01636(.a(n1426), .b(n1255), .O(n1721));
  andx  g01637(.a(n1426), .b(n1255), .O(n1722));
  orx   g01638(.a(n1722), .b(n1394), .O(n1723));
  andx  g01639(.a(n1723), .b(n1721), .O(n1724));
  andx  g01640(.a(n1724), .b(n1720), .O(n1725));
  orx   g01641(.a(n1725), .b(n1719), .O(n1726));
  andx  g01642(.a(n1383), .b(n255), .O(n1727));
  andx  g01643(.a(n1408), .b(n1403), .O(n1728));
  andx  g01644(.a(n1410), .b(n1404), .O(n1729));
  orx   g01645(.a(n1729), .b(n1728), .O(n1730));
  andx  g01646(.a(n1730), .b(n1398), .O(n1731));
  andx  g01647(.a(n1730), .b(n1246), .O(n1732));
  andx  g01648(.a(n1398), .b(n1246), .O(n1733));
  orx   g01649(.a(n1733), .b(n1732), .O(n1734));
  orx   g01650(.a(n1734), .b(n1731), .O(n1735));
  orx   g01651(.a(n1735), .b(n1727), .O(n1736));
  orx   g01652(.a(n1412), .b(n1400), .O(n1740));
  orx   g01653(.a(n1412), .b(n1397), .O(n1741));
  orx   g01654(.a(n1400), .b(n1397), .O(n1742));
  andx  g01655(.a(n1742), .b(n1741), .O(n1743));
  andx  g01656(.a(n1743), .b(n1740), .O(n1744));
  orx   g01657(.a(n1744), .b(n1393), .O(n1745));
  andx  g01658(.a(n1745), .b(n1736), .O(n1746));
  orx   g01659(.a(n1251), .b(n481), .O(n1747));
  orx   g01660(.a(n1747), .b(n1411), .O(n1748));
  invx  g01661(.a(n1411), .O(n1749));
  andx  g01662(.a(n1238), .b(n499), .O(n1750));
  orx   g01663(.a(n1750), .b(n1749), .O(n1751));
  andx  g01664(.a(n1751), .b(n1748), .O(n1752));
  andx  g01665(.a(n914), .b(n554), .O(n1753));
  invx  g01666(.a(n1753), .O(n1754));
  orx   g01667(.a(n1407), .b(n477), .O(n1755));
  andx  g01668(.a(n1755), .b(n1754), .O(n1756));
  andx  g01669(.a(n1084), .b(n488), .O(n1757));
  andx  g01670(.a(n1757), .b(n1753), .O(n1758));
  orx   g01671(.a(n1758), .b(n1756), .O(n1759));
  andx  g01672(.a(n1759), .b(n1752), .O(n1760));
  andx  g01673(.a(n1750), .b(n1749), .O(n1761));
  andx  g01674(.a(n1747), .b(n1411), .O(n1762));
  orx   g01675(.a(n1762), .b(n1761), .O(n1763));
  andx  g01676(.a(n2380), .b(n1763), .O(n1765));
  orx   g01677(.a(n1765), .b(n1760), .O(n1766));
  orx   g01678(.a(n1766), .b(n1746), .O(n1767));
  orx   g01679(.a(n1393), .b(n254), .O(n1768));
  andx  g01680(.a(n1744), .b(n1768), .O(n1769));
  andx  g01681(.a(n1735), .b(n1383), .O(n1770));
  orx   g01682(.a(n1770), .b(n1769), .O(n1771));
  orx   g01683(.a(n2380), .b(n1763), .O(n1772));
  orx   g01684(.a(n1759), .b(n1752), .O(n1773));
  andx  g01685(.a(n1773), .b(n1772), .O(n1774));
  orx   g01686(.a(n1774), .b(n1771), .O(n1775));
  andx  g01687(.a(n1775), .b(n1767), .O(n1776));
  orx   g01688(.a(n1776), .b(n1726), .O(n1777));
  orx   g01689(.a(n1724), .b(n1720), .O(n1778));
  orx   g01690(.a(n1718), .b(n1714), .O(n1779));
  andx  g01691(.a(n1779), .b(n1778), .O(n1780));
  andx  g01692(.a(n1774), .b(n1771), .O(n1781));
  andx  g01693(.a(n1766), .b(n1746), .O(n1782));
  orx   g01694(.a(n1782), .b(n1781), .O(n1783));
  orx   g01695(.a(n1783), .b(n1780), .O(n1784));
  andx  g01696(.a(n1784), .b(n1777), .O(n1785));
  andx  g01697(.a(n1785), .b(n1713), .O(n1786));
  invx  g01698(.a(n1786), .O(n1787));
  orx   g01699(.a(n1785), .b(n1713), .O(n1788));
  andx  g01700(.a(n1788), .b(n1787), .O(n1789));
  invx  g01701(.a(n1789), .O(n1790));
  orx   g01702(.a(n1557), .b(n1554), .O(n1791));
  orx   g01703(.a(n1552), .b(n1429), .O(n1792));
  andx  g01704(.a(n1792), .b(n1791), .O(n1793));
  andx  g01705(.a(n1559), .b(n836), .O(n1794));
  andx  g01706(.a(n1238), .b(n836), .O(n1795));
  andx  g01707(.a(n1795), .b(n1084), .O(n1796));
  andx  g01708(.a(n1084), .b(n836), .O(n1797));
  andx  g01709(.a(n1797), .b(n914), .O(n1798));
  orx   g01710(.a(n1798), .b(n1796), .O(n1799));
  andx  g01711(.a(n1799), .b(n1383), .O(n1800));
  andx  g01712(.a(n1238), .b(n835), .O(n1801));
  andx  g01713(.a(n1383), .b(n836), .O(n1802));
  orx   g01714(.a(n1802), .b(n1799), .O(n1803));
  andx  g01715(.a(n1803), .b(n1801), .O(n1804));
  orx   g01716(.a(n1804), .b(n1800), .O(n1805));
  andx  g01717(.a(n1805), .b(n1794), .O(n1806));
  invx  g01718(.a(n1806), .O(n1807));
  invx  g01719(.a(n1794), .O(n1808));
  invx  g01720(.a(n1805), .O(n1809));
  andx  g01721(.a(n1809), .b(n1808), .O(n1810));
  orx   g01722(.a(n1810), .b(n1393), .O(n1811));
  andx  g01723(.a(n1811), .b(n1807), .O(n1812));
  andx  g01724(.a(n1698), .b(n836), .O(n1813));
  invx  g01725(.a(n1813), .O(n1814));
  andx  g01726(.a(n1814), .b(n1812), .O(n1815));
  invx  g01727(.a(n1812), .O(n1816));
  andx  g01728(.a(n1813), .b(n1816), .O(n1817));
  orx   g01729(.a(n1817), .b(n1815), .O(n1818));
  invx  g01730(.a(n1818), .O(n1819));
  andx  g01731(.a(n1819), .b(n1793), .O(n1820));
  andx  g01732(.a(n1818), .b(n1559), .O(n1821));
  orx   g01733(.a(n1821), .b(n1820), .O(n1822));
  andx  g01734(.a(n1692), .b(n1594), .O(n1823));
  invx  g01735(.a(n1823), .O(n1824));
  andx  g01736(.a(n1680), .b(n1556), .O(n1825));
  orx   g01737(.a(n1825), .b(n1681), .O(n1826));
  orx   g01738(.a(n1826), .b(n1683), .O(n1827));
  andx  g01739(.a(n1653), .b(n1642), .O(n1828));
  orx   g01740(.a(n1828), .b(n1659), .O(n1829));
  invx  g01741(.a(n1829), .O(n1830));
  andx  g01742(.a(n1830), .b(n488), .O(n1831));
  invx  g01743(.a(n1831), .O(n1832));
  andx  g01744(.a(n836), .b(n338), .O(n1833));
  invx  g01745(.a(n1833), .O(n1834));
  andx  g01746(.a(n1616), .b(n1613), .O(n1835));
  invx  g01747(.a(n1835), .O(n1836));
  andx  g01748(.a(n1836), .b(n1614), .O(n1837));
  andx  g01749(.a(n1837), .b(n467), .O(n1841));
  invx  g01750(.a(n1841), .O(n1842));
  andx  g01751(.a(n1842), .b(n1836), .O(n1843));
  invx  g01752(.a(n1843), .O(n1844));
  andx  g01753(.a(n1844), .b(n1834), .O(n1845));
  andx  g01754(.a(n1843), .b(n1833), .O(n1846));
  orx   g01755(.a(n1846), .b(n1845), .O(n1847));
  invx  g01756(.a(n1629), .O(n1848));
  andx  g01757(.a(n1848), .b(n1622), .O(n1849));
  andx  g01758(.a(n1629), .b(n1621), .O(n1850));
  invx  g01759(.a(n1850), .O(n1851));
  andx  g01760(.a(n1851), .b(n1623), .O(n1852));
  orx   g01761(.a(n1852), .b(n1849), .O(n1853));
  andx  g01762(.a(n559), .b(n299), .O(n1854));
  orx   g01763(.a(n1854), .b(n1853), .O(n1855));
  andx  g01764(.a(n1855), .b(n1847), .O(n1856));
  invx  g01765(.a(n1856), .O(n1857));
  orx   g01766(.a(n1855), .b(n1847), .O(n1858));
  andx  g01767(.a(n1858), .b(n1857), .O(n1859));
  invx  g01768(.a(n1859), .O(n1860));
  andx  g01769(.a(n1637), .b(n1493), .O(n1861));
  invx  g01770(.a(n1861), .O(n1862));
  andx  g01771(.a(n1640), .b(n1479), .O(n1863));
  orx   g01772(.a(n1863), .b(n1603), .O(n1864));
  andx  g01773(.a(n1864), .b(n1862), .O(n1865));
  andx  g01774(.a(n827), .b(n554), .O(n1866));
  invx  g01775(.a(n1866), .O(n1867));
  andx  g01776(.a(n1867), .b(n1865), .O(n1868));
  invx  g01777(.a(n1865), .O(n1869));
  andx  g01778(.a(n1866), .b(n1869), .O(n1870));
  orx   g01779(.a(n1870), .b(n1868), .O(n1871));
  orx   g01780(.a(n1871), .b(n1860), .O(n1872));
  andx  g01781(.a(n1871), .b(n1860), .O(n1873));
  invx  g01782(.a(n1873), .O(n1874));
  andx  g01783(.a(n1874), .b(n1872), .O(n1875));
  andx  g01784(.a(n1875), .b(n1832), .O(n1876));
  invx  g01785(.a(n1872), .O(n1877));
  orx   g01786(.a(n1873), .b(n1877), .O(n1878));
  andx  g01787(.a(n1878), .b(n1831), .O(n1879));
  orx   g01788(.a(n1879), .b(n1876), .O(n1880));
  andx  g01789(.a(n1664), .b(n499), .O(n1881));
  orx   g01790(.a(n1881), .b(n1597), .O(n1882));
  andx  g01791(.a(n1882), .b(n1880), .O(n1883));
  orx   g01792(.a(n1878), .b(n1831), .O(n1884));
  orx   g01793(.a(n1875), .b(n1832), .O(n1885));
  andx  g01794(.a(n1885), .b(n1884), .O(n1886));
  invx  g01795(.a(n1882), .O(n1887));
  andx  g01796(.a(n1887), .b(n1886), .O(n1888));
  orx   g01797(.a(n1888), .b(n1883), .O(n1889));
  andx  g01798(.a(n1889), .b(n1827), .O(n1890));
  invx  g01799(.a(n1827), .O(n1891));
  orx   g01800(.a(n1887), .b(n1886), .O(n1892));
  orx   g01801(.a(n1882), .b(n1880), .O(n1893));
  andx  g01802(.a(n1893), .b(n1892), .O(n1894));
  andx  g01803(.a(n1894), .b(n1891), .O(n1895));
  orx   g01804(.a(n1895), .b(n1890), .O(n1896));
  andx  g01805(.a(n1896), .b(n1824), .O(n1897));
  orx   g01806(.a(n1894), .b(n1891), .O(n1898));
  orx   g01807(.a(n1889), .b(n1827), .O(n1899));
  andx  g01808(.a(n1899), .b(n1898), .O(n1900));
  andx  g01809(.a(n1900), .b(n1823), .O(n1901));
  orx   g01810(.a(n1901), .b(n1897), .O(n1902));
  andx  g01811(.a(n1902), .b(n605), .O(n1903));
  invx  g01812(.a(n1903), .O(n1904));
  andx  g01813(.a(n1809), .b(n1794), .O(n1905));
  andx  g01814(.a(n1805), .b(n1808), .O(n1906));
  orx   g01815(.a(n1906), .b(n1905), .O(n1907));
  andx  g01816(.a(n1907), .b(n1383), .O(n1908));
  invx  g01817(.a(n1908), .O(n1909));
  orx   g01818(.a(n1907), .b(n1383), .O(n1910));
  andx  g01819(.a(n1910), .b(n1909), .O(n1911));
  invx  g01820(.a(n1800), .O(n1912));
  andx  g01821(.a(n1803), .b(n1912), .O(n1913));
  invx  g01822(.a(n1913), .O(n1914));
  andx  g01823(.a(n1914), .b(n1801), .O(n1915));
  invx  g01824(.a(n1915), .O(n1916));
  orx   g01825(.a(n1914), .b(n1801), .O(n1917));
  andx  g01826(.a(n1917), .b(n1916), .O(n1918));
  invx  g01827(.a(n1918), .O(n1919));
  andx  g01828(.a(n1797), .b(n1079), .O(n1920));
  invx  g01829(.a(n1920), .O(n1921));
  orx   g01830(.a(n1797), .b(n1079), .O(n1922));
  andx  g01831(.a(n1922), .b(n1921), .O(n1923));
  invx  g01832(.a(n1923), .O(n1924));
  andx  g01833(.a(n1238), .b(n605), .O(n1925));
  andx  g01834(.a(n1925), .b(n1924), .O(n1926));
  andx  g01835(.a(n914), .b(n836), .O(n1927));
  andx  g01836(.a(n1084), .b(n605), .O(n1928));
  andx  g01837(.a(n1928), .b(n1927), .O(n1929));
  andx  g01838(.a(n1929), .b(n1925), .O(n1930));
  orx   g01839(.a(n1930), .b(n1926), .O(n1931));
  andx  g01840(.a(n1931), .b(n1383), .O(n1932));
  orx   g01841(.a(n1798), .b(n1795), .O(n1933));
  andx  g01842(.a(n1798), .b(n1795), .O(n1934));
  invx  g01843(.a(n1934), .O(n1935));
  andx  g01844(.a(n1935), .b(n1933), .O(n1936));
  invx  g01845(.a(n1936), .O(n1937));
  andx  g01846(.a(n1937), .b(n1407), .O(n1938));
  andx  g01847(.a(n1936), .b(n1084), .O(n1939));
  orx   g01848(.a(n1939), .b(n1938), .O(n1940));
  invx  g01849(.a(n1940), .O(n1941));
  andx  g01850(.a(n1383), .b(n605), .O(n1942));
  orx   g01851(.a(n1942), .b(n1931), .O(n1943));
  andx  g01852(.a(n1943), .b(n1941), .O(n1944));
  orx   g01853(.a(n1944), .b(n1932), .O(n1945));
  andx  g01854(.a(n1945), .b(n1919), .O(n1946));
  invx  g01855(.a(n1946), .O(n1947));
  andx  g01856(.a(n1559), .b(n605), .O(n1948));
  invx  g01857(.a(n1948), .O(n1949));
  invx  g01858(.a(n1945), .O(n1950));
  andx  g01859(.a(n1950), .b(n1918), .O(n1951));
  orx   g01860(.a(n1951), .b(n1949), .O(n1952));
  andx  g01861(.a(n1952), .b(n1947), .O(n1953));
  invx  g01862(.a(n1953), .O(n1954));
  andx  g01863(.a(n1954), .b(n1911), .O(n1955));
  orx   g01864(.a(n1954), .b(n1911), .O(n1956));
  andx  g01865(.a(n1698), .b(n605), .O(n1957));
  andx  g01866(.a(n1957), .b(n1956), .O(n1958));
  orx   g01867(.a(n1958), .b(n1955), .O(n1959));
  andx  g01868(.a(n1959), .b(n1904), .O(n1960));
  invx  g01869(.a(n1960), .O(n1961));
  orx   g01870(.a(n1959), .b(n1904), .O(n1962));
  andx  g01871(.a(n1962), .b(n1961), .O(n1963));
  orx   g01872(.a(n1963), .b(n1822), .O(n1964));
  invx  g01873(.a(n1964), .O(n1965));
  andx  g01874(.a(n1963), .b(n1822), .O(n1966));
  orx   g01875(.a(n1966), .b(n1965), .O(n1967));
  invx  g01876(.a(n1957), .O(n1968));
  andx  g01877(.a(n1968), .b(n1953), .O(n1969));
  andx  g01878(.a(n1957), .b(n1954), .O(n1970));
  orx   g01879(.a(n1970), .b(n1969), .O(n1971));
  orx   g01880(.a(n1971), .b(n1911), .O(n1972));
  invx  g01881(.a(n1972), .O(n1973));
  andx  g01882(.a(n1971), .b(n1911), .O(n1974));
  orx   g01883(.a(n1974), .b(n1973), .O(n1975));
  orx   g01884(.a(n1948), .b(n1945), .O(n1976));
  andx  g01885(.a(n1948), .b(n1945), .O(n1977));
  invx  g01886(.a(n1977), .O(n1978));
  andx  g01887(.a(n1978), .b(n1976), .O(n1979));
  andx  g01888(.a(n1979), .b(n1918), .O(n1980));
  invx  g01889(.a(n1976), .O(n1981));
  orx   g01890(.a(n1977), .b(n1981), .O(n1982));
  andx  g01891(.a(n1982), .b(n1919), .O(n1983));
  orx   g01892(.a(n1983), .b(n1980), .O(n1984));
  invx  g01893(.a(n1932), .O(n1985));
  andx  g01894(.a(n1943), .b(n1985), .O(n1986));
  invx  g01895(.a(n1986), .O(n1987));
  andx  g01896(.a(n1987), .b(n1941), .O(n1988));
  andx  g01897(.a(n1986), .b(n1940), .O(n1989));
  orx   g01898(.a(n1989), .b(n1988), .O(n1990));
  andx  g01899(.a(n1238), .b(n554), .O(n1991));
  invx  g01900(.a(n1927), .O(n1992));
  orx   g01901(.a(n1928), .b(n1992), .O(n1993));
  invx  g01902(.a(n1993), .O(n1994));
  andx  g01903(.a(n1928), .b(n1992), .O(n1995));
  orx   g01904(.a(n1995), .b(n1994), .O(n1996));
  andx  g01905(.a(n1996), .b(n1991), .O(n1997));
  andx  g01906(.a(n914), .b(n605), .O(n1998));
  andx  g01907(.a(n1084), .b(n554), .O(n1999));
  andx  g01908(.a(n1999), .b(n1998), .O(n2000));
  andx  g01909(.a(n2000), .b(n1991), .O(n2001));
  andx  g01910(.a(n2000), .b(n1996), .O(n2002));
  orx   g01911(.a(n2002), .b(n2001), .O(n2003));
  orx   g01912(.a(n2003), .b(n1997), .O(n2004));
  andx  g01913(.a(n2004), .b(n1383), .O(n2005));
  invx  g01914(.a(n1929), .O(n2006));
  andx  g01915(.a(n2006), .b(n1925), .O(n2007));
  invx  g01916(.a(n2007), .O(n2008));
  orx   g01917(.a(n2006), .b(n1925), .O(n2009));
  andx  g01918(.a(n2009), .b(n2008), .O(n2010));
  andx  g01919(.a(n2010), .b(n1924), .O(n2011));
  invx  g01920(.a(n2009), .O(n2012));
  orx   g01921(.a(n2012), .b(n2007), .O(n2013));
  andx  g01922(.a(n2013), .b(n1923), .O(n2014));
  orx   g01923(.a(n2014), .b(n2011), .O(n2015));
  andx  g01924(.a(n1383), .b(n554), .O(n2016));
  orx   g01925(.a(n2016), .b(n2004), .O(n2017));
  andx  g01926(.a(n2017), .b(n2015), .O(n2018));
  orx   g01927(.a(n2018), .b(n2005), .O(n2019));
  andx  g01928(.a(n2019), .b(n1990), .O(n2020));
  andx  g01929(.a(n1559), .b(n554), .O(n2021));
  orx   g01930(.a(n2019), .b(n1990), .O(n2022));
  andx  g01931(.a(n2022), .b(n2021), .O(n2023));
  orx   g01932(.a(n2023), .b(n2020), .O(n2024));
  andx  g01933(.a(n2024), .b(n1984), .O(n2025));
  orx   g01934(.a(n2024), .b(n1984), .O(n2026));
  andx  g01935(.a(n1698), .b(n554), .O(n2027));
  andx  g01936(.a(n2027), .b(n2026), .O(n2028));
  orx   g01937(.a(n2028), .b(n2025), .O(n2029));
  andx  g01938(.a(n2029), .b(n1975), .O(n2030));
  invx  g01939(.a(n2030), .O(n2031));
  andx  g01940(.a(n1902), .b(n554), .O(n2032));
  invx  g01941(.a(n2032), .O(n2033));
  invx  g01942(.a(n1974), .O(n2034));
  andx  g01943(.a(n2034), .b(n1972), .O(n2035));
  invx  g01944(.a(n2025), .O(n2036));
  orx   g01945(.a(n1982), .b(n1919), .O(n2037));
  orx   g01946(.a(n1979), .b(n1918), .O(n2038));
  andx  g01947(.a(n2038), .b(n2037), .O(n2039));
  invx  g01948(.a(n2024), .O(n2040));
  andx  g01949(.a(n2040), .b(n2039), .O(n2041));
  invx  g01950(.a(n2027), .O(n2042));
  orx   g01951(.a(n2042), .b(n2041), .O(n2043));
  andx  g01952(.a(n2043), .b(n2036), .O(n2044));
  andx  g01953(.a(n2044), .b(n2035), .O(n2045));
  orx   g01954(.a(n2045), .b(n2033), .O(n2046));
  andx  g01955(.a(n2046), .b(n2031), .O(n2047));
  andx  g01956(.a(n1896), .b(n1823), .O(n2048));
  invx  g01957(.a(n2048), .O(n2049));
  andx  g01958(.a(n1882), .b(n1886), .O(n2053));
  andx  g01959(.a(n1878), .b(n488), .O(n2054));
  orx   g01960(.a(n2054), .b(n1829), .O(n2055));
  andx  g01961(.a(n836), .b(n299), .O(n2056));
  invx  g01962(.a(n2056), .O(n2057));
  andx  g01963(.a(n1842), .b(n1833), .O(n2058));
  orx   g01964(.a(n2058), .b(n1835), .O(n2059));
  invx  g01965(.a(n2059), .O(n2060));
  andx  g01966(.a(n2060), .b(n551), .O(n2061));
  invx  g01967(.a(n2061), .O(n2062));
  invx  g01968(.a(n2058), .O(n2064));
  andx  g01969(.a(n2064), .b(n2062), .O(n2065));
  invx  g01970(.a(n2065), .O(n2066));
  andx  g01971(.a(n2066), .b(n2057), .O(n2067));
  andx  g01972(.a(n2065), .b(n2056), .O(n2068));
  orx   g01973(.a(n2068), .b(n2067), .O(n2069));
  invx  g01974(.a(n1847), .O(n2070));
  andx  g01975(.a(n1853), .b(n2070), .O(n2071));
  andx  g01976(.a(n2071), .b(n827), .O(n2072));
  invx  g01977(.a(n2072), .O(n2073));
  andx  g01978(.a(n827), .b(n605), .O(n2074));
  orx   g01979(.a(n2074), .b(n2071), .O(n2075));
  andx  g01980(.a(n2075), .b(n2073), .O(n2076));
  invx  g01981(.a(n2076), .O(n2077));
  andx  g01982(.a(n2077), .b(n2069), .O(n2078));
  invx  g01983(.a(n2069), .O(n2079));
  andx  g01984(.a(n2076), .b(n2079), .O(n2080));
  orx   g01985(.a(n2080), .b(n2078), .O(n2081));
  andx  g01986(.a(n1869), .b(n1860), .O(n2082));
  invx  g01987(.a(n2082), .O(n2083));
  andx  g01988(.a(n1865), .b(n1859), .O(n2084));
  orx   g01989(.a(n2084), .b(n1867), .O(n2085));
  andx  g01990(.a(n2085), .b(n2083), .O(n2086));
  andx  g01991(.a(n2086), .b(n554), .O(n2087));
  invx  g01992(.a(n2087), .O(n2088));
  andx  g01993(.a(n2088), .b(n2081), .O(n2089));
  invx  g01994(.a(n2081), .O(n2090));
  andx  g01995(.a(n2087), .b(n2090), .O(n2091));
  orx   g01996(.a(n2091), .b(n2089), .O(n2092));
  invx  g01997(.a(n2092), .O(n2093));
  andx  g01998(.a(n2093), .b(n2055), .O(n2094));
  orx   g01999(.a(n2093), .b(n2055), .O(n2095));
  invx  g02000(.a(n2095), .O(n2096));
  orx   g02001(.a(n2096), .b(n2094), .O(n2097));
  orx   g02002(.a(n2097), .b(n2053), .O(n2098));
  orx   g02003(.a(n2098), .b(n1890), .O(n2099));
  invx  g02004(.a(n2053), .O(n2100));
  invx  g02005(.a(n2094), .O(n2101));
  andx  g02006(.a(n2095), .b(n2101), .O(n2102));
  orx   g02007(.a(n2102), .b(n2100), .O(n2103));
  orx   g02008(.a(n2102), .b(n1898), .O(n2105));
  andx  g02009(.a(n2105), .b(n2103), .O(n2106));
  andx  g02010(.a(n2106), .b(n2099), .O(n2107));
  andx  g02011(.a(n2107), .b(n2049), .O(n2108));
  andx  g02012(.a(n2102), .b(n2100), .O(n2109));
  andx  g02013(.a(n2109), .b(n1898), .O(n2110));
  andx  g02014(.a(n2097), .b(n2053), .O(n2111));
  andx  g02015(.a(n2097), .b(n1890), .O(n2112));
  orx   g02016(.a(n2112), .b(n2111), .O(n2113));
  orx   g02017(.a(n2113), .b(n2110), .O(n2114));
  andx  g02018(.a(n2114), .b(n2048), .O(n2115));
  orx   g02019(.a(n2115), .b(n2108), .O(n2116));
  andx  g02020(.a(n2116), .b(n554), .O(n2117));
  orx   g02021(.a(n2117), .b(n2047), .O(n2118));
  orx   g02022(.a(n2029), .b(n1975), .O(n2119));
  andx  g02023(.a(n2119), .b(n2032), .O(n2120));
  orx   g02024(.a(n2120), .b(n2030), .O(n2121));
  invx  g02025(.a(n2117), .O(n2122));
  orx   g02026(.a(n2122), .b(n2121), .O(n2123));
  andx  g02027(.a(n2123), .b(n2118), .O(n2124));
  orx   g02028(.a(n2124), .b(n1967), .O(n2125));
  invx  g02029(.a(n1966), .O(n2126));
  andx  g02030(.a(n2126), .b(n1964), .O(n2127));
  andx  g02031(.a(n2122), .b(n2121), .O(n2128));
  andx  g02032(.a(n2117), .b(n2047), .O(n2129));
  orx   g02033(.a(n2129), .b(n2128), .O(n2130));
  orx   g02034(.a(n2130), .b(n2127), .O(n2131));
  andx  g02035(.a(n2131), .b(n2125), .O(n2132));
  andx  g02036(.a(n2107), .b(n2048), .O(n2133));
  invx  g02037(.a(n2133), .O(n2134));
  andx  g02038(.a(n2100), .b(n1898), .O(n2135));
  orx   g02039(.a(n2135), .b(n2097), .O(n2136));
  andx  g02040(.a(n2062), .b(n2056), .O(n2137));
  orx   g02041(.a(n2137), .b(n2058), .O(n2138));
  invx  g02042(.a(n2138), .O(n2139));
  andx  g02043(.a(n827), .b(n610), .O(n2140));
  invx  g02044(.a(n2140), .O(n2141));
  andx  g02045(.a(n2141), .b(n2139), .O(n2142));
  invx  g02046(.a(n2142), .O(n2143));
  andx  g02047(.a(n2143), .b(n602), .O(n2144));
  andx  g02048(.a(n2142), .b(n299), .O(n2145));
  orx   g02049(.a(n2145), .b(n2144), .O(n2146));
  invx  g02050(.a(n2146), .O(n2147));
  andx  g02051(.a(n2075), .b(n2079), .O(n2148));
  orx   g02052(.a(n2148), .b(n2072), .O(n2149));
  invx  g02053(.a(n2149), .O(n2150));
  andx  g02054(.a(n2150), .b(n605), .O(n2151));
  invx  g02055(.a(n2151), .O(n2152));
  andx  g02056(.a(n2152), .b(n2147), .O(n2153));
  orx   g02057(.a(n2439), .b(n2153), .O(n2155));
  andx  g02058(.a(n2090), .b(n554), .O(n2156));
  invx  g02059(.a(n2156), .O(n2157));
  andx  g02060(.a(n2157), .b(n2086), .O(n2158));
  invx  g02061(.a(n2155), .O(n2161));
  andx  g02062(.a(n2158), .b(n2161), .O(n2162));
  invx  g02063(.a(n2162), .O(n2164));
  orx   g02064(.a(n2094), .b(n2164), .O(n2167));
  andx  g02065(.a(n2167), .b(n2136), .O(n2168));
  orx   g02066(.a(n2167), .b(n2136), .O(n2169));
  orx   g02067(.a(n2452), .b(n2168), .O(n2171));
  andx  g02068(.a(n2171), .b(n2134), .O(n2172));
  invx  g02069(.a(n2168), .O(n2173));
  andx  g02070(.a(n2169), .b(n2173), .O(n2174));
  andx  g02071(.a(n2174), .b(n2133), .O(n2175));
  orx   g02072(.a(n2175), .b(n2172), .O(n2176));
  andx  g02073(.a(n2033), .b(n2029), .O(n2177));
  andx  g02074(.a(n2032), .b(n2044), .O(n2178));
  orx   g02075(.a(n2178), .b(n2177), .O(n2179));
  andx  g02076(.a(n2179), .b(n2035), .O(n2180));
  orx   g02077(.a(n2032), .b(n2044), .O(n2181));
  orx   g02078(.a(n2033), .b(n2029), .O(n2182));
  andx  g02079(.a(n2182), .b(n2181), .O(n2183));
  andx  g02080(.a(n2183), .b(n1975), .O(n2184));
  orx   g02081(.a(n2184), .b(n2180), .O(n2185));
  orx   g02082(.a(n2027), .b(n2024), .O(n2186));
  andx  g02083(.a(n2027), .b(n2024), .O(n2187));
  invx  g02084(.a(n2187), .O(n2188));
  andx  g02085(.a(n2188), .b(n2186), .O(n2189));
  andx  g02086(.a(n2189), .b(n2039), .O(n2190));
  invx  g02087(.a(n2186), .O(n2191));
  orx   g02088(.a(n2187), .b(n2191), .O(n2192));
  andx  g02089(.a(n2192), .b(n1984), .O(n2193));
  orx   g02090(.a(n2193), .b(n2190), .O(n2194));
  invx  g02091(.a(n1990), .O(n2195));
  orx   g02092(.a(n2021), .b(n2019), .O(n2196));
  invx  g02093(.a(n2196), .O(n2197));
  andx  g02094(.a(n2021), .b(n2019), .O(n2198));
  orx   g02095(.a(n2198), .b(n2197), .O(n2199));
  orx   g02096(.a(n2199), .b(n2195), .O(n2200));
  invx  g02097(.a(n2198), .O(n2201));
  andx  g02098(.a(n2201), .b(n2196), .O(n2202));
  orx   g02099(.a(n2202), .b(n1990), .O(n2203));
  andx  g02100(.a(n2203), .b(n2200), .O(n2204));
  orx   g02101(.a(n2013), .b(n1923), .O(n2205));
  orx   g02102(.a(n2010), .b(n1924), .O(n2206));
  andx  g02103(.a(n2206), .b(n2205), .O(n2207));
  invx  g02104(.a(n1997), .O(n2208));
  orx   g02105(.a(n1251), .b(n560), .O(n2209));
  invx  g02106(.a(n2000), .O(n2210));
  orx   g02107(.a(n2210), .b(n2209), .O(n2211));
  invx  g02108(.a(n1995), .O(n2212));
  andx  g02109(.a(n2212), .b(n1993), .O(n2213));
  orx   g02110(.a(n2210), .b(n2213), .O(n2214));
  andx  g02111(.a(n2214), .b(n2211), .O(n2215));
  andx  g02112(.a(n2215), .b(n2208), .O(n2216));
  orx   g02113(.a(n2216), .b(n1393), .O(n2217));
  andx  g02114(.a(n2017), .b(n2217), .O(n2218));
  orx   g02115(.a(n2218), .b(n2207), .O(n2219));
  orx   g02116(.a(n1393), .b(n560), .O(n2220));
  andx  g02117(.a(n2220), .b(n2216), .O(n2221));
  orx   g02118(.a(n2221), .b(n2005), .O(n2222));
  orx   g02119(.a(n2222), .b(n2015), .O(n2223));
  andx  g02120(.a(n2223), .b(n2219), .O(n2224));
  orx   g02121(.a(n1393), .b(n477), .O(n2225));
  andx  g02122(.a(n1238), .b(n488), .O(n2226));
  andx  g02123(.a(n2226), .b(n1758), .O(n2227));
  invx  g02124(.a(n2227), .O(n2228));
  invx  g02125(.a(n1758), .O(n2229));
  invx  g02126(.a(n1998), .O(n2230));
  orx   g02127(.a(n1999), .b(n2230), .O(n2231));
  andx  g02128(.a(n1999), .b(n2230), .O(n2232));
  invx  g02129(.a(n2232), .O(n2233));
  andx  g02130(.a(n2233), .b(n2231), .O(n2234));
  orx   g02131(.a(n2234), .b(n2229), .O(n2235));
  orx   g02132(.a(n1251), .b(n477), .O(n2236));
  orx   g02133(.a(n2234), .b(n2236), .O(n2237));
  andx  g02134(.a(n2237), .b(n2235), .O(n2238));
  andx  g02135(.a(n2238), .b(n2228), .O(n2239));
  andx  g02136(.a(n2239), .b(n2225), .O(n2240));
  andx  g02137(.a(n2210), .b(n1991), .O(n2241));
  andx  g02138(.a(n2000), .b(n2209), .O(n2242));
  orx   g02139(.a(n2242), .b(n2241), .O(n2243));
  orx   g02140(.a(n1996), .b(n2243), .O(n2248));
  invx  g02141(.a(n2248), .O(n2249));
  andx  g02142(.a(n1996), .b(n2243), .O(n2250));
  orx   g02143(.a(n2250), .b(n2249), .O(n2251));
  orx   g02144(.a(n2251), .b(n2240), .O(n2252));
  orx   g02145(.a(n2239), .b(n1393), .O(n2253));
  andx  g02146(.a(n2253), .b(n2252), .O(n2254));
  andx  g02147(.a(n2254), .b(n2224), .O(n2255));
  invx  g02148(.a(n2255), .O(n2256));
  andx  g02149(.a(n2222), .b(n2015), .O(n2257));
  andx  g02150(.a(n2218), .b(n2207), .O(n2258));
  orx   g02151(.a(n2258), .b(n2257), .O(n2259));
  andx  g02152(.a(n1559), .b(n488), .O(n2260));
  orx   g02153(.a(n2260), .b(n2259), .O(n2261));
  andx  g02154(.a(n1383), .b(n488), .O(n2262));
  invx  g02155(.a(n2231), .O(n2263));
  orx   g02156(.a(n2232), .b(n2263), .O(n2264));
  andx  g02157(.a(n2264), .b(n1758), .O(n2265));
  andx  g02158(.a(n2264), .b(n2226), .O(n2266));
  orx   g02159(.a(n2266), .b(n2265), .O(n2267));
  orx   g02160(.a(n2267), .b(n2227), .O(n2268));
  orx   g02161(.a(n2268), .b(n2262), .O(n2269));
  invx  g02162(.a(n2250), .O(n2270));
  andx  g02163(.a(n2270), .b(n2248), .O(n2271));
  andx  g02164(.a(n2271), .b(n2269), .O(n2272));
  andx  g02165(.a(n2268), .b(n1383), .O(n2273));
  orx   g02166(.a(n2273), .b(n2272), .O(n2274));
  orx   g02167(.a(n2260), .b(n2274), .O(n2275));
  andx  g02168(.a(n2275), .b(n2261), .O(n2276));
  andx  g02169(.a(n2276), .b(n2256), .O(n2277));
  andx  g02170(.a(n2277), .b(n2204), .O(n2278));
  orx   g02171(.a(n2277), .b(n2204), .O(n2279));
  andx  g02172(.a(n1698), .b(n488), .O(n2280));
  andx  g02173(.a(n2280), .b(n2279), .O(n2281));
  orx   g02174(.a(n2281), .b(n2278), .O(n2282));
  andx  g02175(.a(n2282), .b(n2194), .O(n2283));
  andx  g02176(.a(n1902), .b(n488), .O(n2284));
  orx   g02177(.a(n2282), .b(n2194), .O(n2285));
  andx  g02178(.a(n2285), .b(n2284), .O(n2286));
  orx   g02179(.a(n2286), .b(n2283), .O(n2287));
  andx  g02180(.a(n2287), .b(n2185), .O(n2288));
  orx   g02181(.a(n2287), .b(n2185), .O(n2289));
  andx  g02182(.a(n2116), .b(n488), .O(n2290));
  andx  g02183(.a(n2290), .b(n2289), .O(n2291));
  orx   g02184(.a(n2291), .b(n2288), .O(n2292));
  andx  g02185(.a(n2292), .b(n2176), .O(n2293));
  invx  g02186(.a(n2288), .O(n2294));
  orx   g02187(.a(n2183), .b(n1975), .O(n2295));
  orx   g02188(.a(n2179), .b(n2035), .O(n2296));
  andx  g02189(.a(n2296), .b(n2295), .O(n2297));
  invx  g02190(.a(n2283), .O(n2298));
  invx  g02191(.a(n2284), .O(n2299));
  orx   g02192(.a(n2192), .b(n1984), .O(n2300));
  orx   g02193(.a(n2189), .b(n2039), .O(n2301));
  andx  g02194(.a(n2301), .b(n2300), .O(n2302));
  invx  g02195(.a(n2278), .O(n2303));
  andx  g02196(.a(n2202), .b(n1990), .O(n2304));
  andx  g02197(.a(n2199), .b(n2195), .O(n2305));
  orx   g02198(.a(n2305), .b(n2304), .O(n2306));
  invx  g02199(.a(n2260), .O(n2307));
  andx  g02200(.a(n2307), .b(n2224), .O(n2308));
  andx  g02201(.a(n2307), .b(n2254), .O(n2309));
  orx   g02202(.a(n2309), .b(n2308), .O(n2310));
  orx   g02203(.a(n2310), .b(n2255), .O(n2311));
  andx  g02204(.a(n2311), .b(n2306), .O(n2312));
  invx  g02205(.a(n2280), .O(n2313));
  orx   g02206(.a(n2313), .b(n2312), .O(n2314));
  andx  g02207(.a(n2314), .b(n2303), .O(n2315));
  andx  g02208(.a(n2315), .b(n2302), .O(n2316));
  orx   g02209(.a(n2316), .b(n2299), .O(n2317));
  andx  g02210(.a(n2317), .b(n2298), .O(n2318));
  andx  g02211(.a(n2318), .b(n2297), .O(n2319));
  invx  g02212(.a(n2290), .O(n2320));
  orx   g02213(.a(n2320), .b(n2319), .O(n2321));
  andx  g02214(.a(n2321), .b(n2294), .O(n2322));
  andx  g02215(.a(n2176), .b(n488), .O(n2323));
  invx  g02216(.a(n2323), .O(n2324));
  andx  g02217(.a(n2324), .b(n2322), .O(n2325));
  orx   g02218(.a(n2325), .b(n2293), .O(n2326));
  andx  g02219(.a(n2326), .b(n2132), .O(n2327));
  andx  g02220(.a(n2130), .b(n2127), .O(n2328));
  andx  g02221(.a(n2124), .b(n1967), .O(n2329));
  orx   g02222(.a(n2329), .b(n2328), .O(n2330));
  orx   g02223(.a(n2174), .b(n2133), .O(n2331));
  orx   g02224(.a(n2171), .b(n2134), .O(n2332));
  andx  g02225(.a(n2332), .b(n2331), .O(n2333));
  orx   g02226(.a(n2322), .b(n2333), .O(n2334));
  orx   g02227(.a(n2323), .b(n2292), .O(n2335));
  andx  g02228(.a(n2335), .b(n2334), .O(n2336));
  andx  g02229(.a(n2336), .b(n2330), .O(n2337));
  orx   g02230(.a(n2337), .b(n2327), .O(n2338));
  orx   g02231(.a(n2290), .b(n2287), .O(n2339));
  orx   g02232(.a(n2320), .b(n2318), .O(n2340));
  andx  g02233(.a(n2340), .b(n2339), .O(n2341));
  andx  g02234(.a(n2341), .b(n2297), .O(n2342));
  andx  g02235(.a(n2320), .b(n2318), .O(n2343));
  andx  g02236(.a(n2290), .b(n2287), .O(n2344));
  orx   g02237(.a(n2344), .b(n2343), .O(n2345));
  andx  g02238(.a(n2345), .b(n2185), .O(n2346));
  orx   g02239(.a(n2346), .b(n2342), .O(n2347));
  orx   g02240(.a(n2284), .b(n2315), .O(n2348));
  orx   g02241(.a(n2299), .b(n2282), .O(n2349));
  andx  g02242(.a(n2349), .b(n2348), .O(n2350));
  orx   g02243(.a(n2350), .b(n2302), .O(n2351));
  andx  g02244(.a(n2299), .b(n2282), .O(n2352));
  andx  g02245(.a(n2284), .b(n2315), .O(n2353));
  orx   g02246(.a(n2353), .b(n2352), .O(n2354));
  orx   g02247(.a(n2354), .b(n2194), .O(n2355));
  andx  g02248(.a(n2355), .b(n2351), .O(n2356));
  andx  g02249(.a(n2280), .b(n2277), .O(n2357));
  andx  g02250(.a(n2313), .b(n2311), .O(n2358));
  orx   g02251(.a(n2358), .b(n2357), .O(n2359));
  orx   g02252(.a(n2359), .b(n2306), .O(n2360));
  orx   g02253(.a(n2313), .b(n2311), .O(n2361));
  orx   g02254(.a(n2280), .b(n2277), .O(n2362));
  andx  g02255(.a(n2362), .b(n2361), .O(n2363));
  orx   g02256(.a(n2363), .b(n2204), .O(n2364));
  andx  g02257(.a(n2364), .b(n2360), .O(n2365));
  andx  g02258(.a(n2260), .b(n2274), .O(n2366));
  orx   g02259(.a(n2366), .b(n2309), .O(n2367));
  orx   g02260(.a(n2367), .b(n2224), .O(n2368));
  orx   g02261(.a(n2307), .b(n2254), .O(n2369));
  andx  g02262(.a(n2369), .b(n2275), .O(n2370));
  orx   g02263(.a(n2370), .b(n2259), .O(n2371));
  andx  g02264(.a(n2371), .b(n2368), .O(n2372));
  andx  g02265(.a(n2253), .b(n2269), .O(n2373));
  orx   g02266(.a(n2373), .b(n2271), .O(n2374));
  orx   g02267(.a(n2273), .b(n2240), .O(n2375));
  orx   g02268(.a(n2375), .b(n2251), .O(n2376));
  andx  g02269(.a(n2376), .b(n2374), .O(n2377));
  andx  g02270(.a(n1755), .b(n1753), .O(n2378));
  andx  g02271(.a(n1757), .b(n1754), .O(n2379));
  orx   g02272(.a(n2379), .b(n2378), .O(n2380));
  andx  g02273(.a(n2380), .b(n1750), .O(n2381));
  andx  g02274(.a(n1750), .b(n1411), .O(n2382));
  andx  g02275(.a(n2380), .b(n1411), .O(n2383));
  orx   g02276(.a(n2383), .b(n2382), .O(n2384));
  orx   g02277(.a(n2384), .b(n2381), .O(n2385));
  andx  g02278(.a(n2385), .b(n1383), .O(n2386));
  andx  g02279(.a(n2226), .b(n2229), .O(n2387));
  andx  g02280(.a(n2236), .b(n1758), .O(n2388));
  orx   g02281(.a(n2388), .b(n2387), .O(n2389));
  orx   g02282(.a(n2264), .b(n2389), .O(n2392));
  orx   g02283(.a(n2236), .b(n1758), .O(n2393));
  orx   g02284(.a(n2226), .b(n2229), .O(n2394));
  andx  g02285(.a(n2394), .b(n2393), .O(n2395));
  orx   g02286(.a(n2234), .b(n2395), .O(n2397));
  andx  g02287(.a(n2397), .b(n2392), .O(n2398));
  andx  g02288(.a(n1383), .b(n499), .O(n2399));
  orx   g02289(.a(n2399), .b(n2385), .O(n2400));
  andx  g02290(.a(n2400), .b(n2398), .O(n2401));
  orx   g02291(.a(n2401), .b(n2386), .O(n2402));
  andx  g02292(.a(n2402), .b(n2377), .O(n2403));
  andx  g02293(.a(n1559), .b(n499), .O(n2404));
  orx   g02294(.a(n2402), .b(n2377), .O(n2405));
  andx  g02295(.a(n2405), .b(n2404), .O(n2406));
  orx   g02296(.a(n2406), .b(n2403), .O(n2407));
  andx  g02297(.a(n2407), .b(n2372), .O(n2408));
  orx   g02298(.a(n2407), .b(n2372), .O(n2409));
  andx  g02299(.a(n1698), .b(n499), .O(n2410));
  andx  g02300(.a(n2410), .b(n2409), .O(n2411));
  orx   g02301(.a(n2411), .b(n2408), .O(n2412));
  andx  g02302(.a(n2412), .b(n2365), .O(n2413));
  andx  g02303(.a(n1902), .b(n499), .O(n2414));
  orx   g02304(.a(n2412), .b(n2365), .O(n2415));
  andx  g02305(.a(n2415), .b(n2414), .O(n2416));
  orx   g02306(.a(n2416), .b(n2413), .O(n2417));
  andx  g02307(.a(n2417), .b(n2356), .O(n2418));
  orx   g02308(.a(n2417), .b(n2356), .O(n2419));
  andx  g02309(.a(n2116), .b(n499), .O(n2420));
  andx  g02310(.a(n2420), .b(n2419), .O(n2421));
  orx   g02311(.a(n2421), .b(n2418), .O(n2422));
  andx  g02312(.a(n2422), .b(n2347), .O(n2423));
  andx  g02313(.a(n2176), .b(n499), .O(n2424));
  orx   g02314(.a(n2422), .b(n2347), .O(n2425));
  andx  g02315(.a(n2425), .b(n2424), .O(n2426));
  orx   g02316(.a(n2426), .b(n2423), .O(n2427));
  andx  g02317(.a(n2171), .b(n2133), .O(n2428));
  invx  g02318(.a(n2428), .O(n2429));
  invx  g02319(.a(n2137), .O(n2432));
  andx  g02320(.a(n2146), .b(n605), .O(n2439));
  invx  g02321(.a(n2136), .O(n2450));
  andx  g02322(.a(n2162), .b(n2450), .O(n2452));
  invx  g02323(.a(n2423), .O(n2465));
  invx  g02324(.a(n2424), .O(n2466));
  orx   g02325(.a(n2345), .b(n2185), .O(n2467));
  orx   g02326(.a(n2341), .b(n2297), .O(n2468));
  andx  g02327(.a(n2468), .b(n2467), .O(n2469));
  invx  g02328(.a(n2418), .O(n2470));
  andx  g02329(.a(n2354), .b(n2194), .O(n2471));
  andx  g02330(.a(n2350), .b(n2302), .O(n2472));
  orx   g02331(.a(n2472), .b(n2471), .O(n2473));
  invx  g02332(.a(n2413), .O(n2474));
  invx  g02333(.a(n2414), .O(n2475));
  andx  g02334(.a(n2363), .b(n2204), .O(n2476));
  andx  g02335(.a(n2359), .b(n2306), .O(n2477));
  orx   g02336(.a(n2477), .b(n2476), .O(n2478));
  invx  g02337(.a(n2408), .O(n2479));
  andx  g02338(.a(n2370), .b(n2259), .O(n2480));
  andx  g02339(.a(n2367), .b(n2224), .O(n2481));
  orx   g02340(.a(n2481), .b(n2480), .O(n2482));
  invx  g02341(.a(n2403), .O(n2483));
  orx   g02342(.a(n1793), .b(n481), .O(n2484));
  andx  g02343(.a(n2375), .b(n2251), .O(n2485));
  andx  g02344(.a(n2373), .b(n2271), .O(n2486));
  orx   g02345(.a(n2486), .b(n2485), .O(n2487));
  orx   g02346(.a(n1759), .b(n1747), .O(n2491));
  orx   g02347(.a(n1747), .b(n1749), .O(n2492));
  orx   g02348(.a(n1759), .b(n1749), .O(n2493));
  andx  g02349(.a(n2493), .b(n2492), .O(n2494));
  andx  g02350(.a(n2494), .b(n2491), .O(n2495));
  orx   g02351(.a(n2495), .b(n1393), .O(n2496));
  andx  g02352(.a(n2234), .b(n2395), .O(n2497));
  andx  g02353(.a(n2264), .b(n2389), .O(n2498));
  orx   g02354(.a(n2498), .b(n2497), .O(n2499));
  orx   g02355(.a(n1393), .b(n481), .O(n2500));
  andx  g02356(.a(n2500), .b(n2495), .O(n2501));
  orx   g02357(.a(n2501), .b(n2499), .O(n2502));
  andx  g02358(.a(n2502), .b(n2496), .O(n2503));
  andx  g02359(.a(n2503), .b(n2487), .O(n2504));
  orx   g02360(.a(n2504), .b(n2484), .O(n2505));
  andx  g02361(.a(n2505), .b(n2483), .O(n2506));
  andx  g02362(.a(n2506), .b(n2482), .O(n2507));
  invx  g02363(.a(n2410), .O(n2508));
  orx   g02364(.a(n2508), .b(n2507), .O(n2509));
  andx  g02365(.a(n2509), .b(n2479), .O(n2510));
  andx  g02366(.a(n2510), .b(n2478), .O(n2511));
  orx   g02367(.a(n2511), .b(n2475), .O(n2512));
  andx  g02368(.a(n2512), .b(n2474), .O(n2513));
  andx  g02369(.a(n2513), .b(n2473), .O(n2514));
  invx  g02370(.a(n2420), .O(n2515));
  orx   g02371(.a(n2515), .b(n2514), .O(n2516));
  andx  g02372(.a(n2516), .b(n2470), .O(n2517));
  andx  g02373(.a(n2517), .b(n2469), .O(n2518));
  orx   g02374(.a(n2518), .b(n2466), .O(n2519));
  andx  g02375(.a(n2519), .b(n2465), .O(n2520));
  andx  g02376(.a(n2520), .b(n499), .O(n2523));
  andx  g02377(.a(n2523), .b(n2338), .O(n2524));
  orx   g02378(.a(n2336), .b(n2330), .O(n2525));
  orx   g02379(.a(n2326), .b(n2132), .O(n2526));
  andx  g02380(.a(n2526), .b(n2525), .O(n2527));
  orx   g02381(.a(n2427), .b(n481), .O(n2530));
  andx  g02382(.a(n2530), .b(n2527), .O(n2531));
  orx   g02383(.a(n2531), .b(n2524), .O(n2532));
  andx  g02384(.a(n2432), .b(n2141), .O(n2535));
  andx  g02385(.a(n2535), .b(n835), .O(n2536));
  invx  g02386(.a(n2536), .O(n2537));
  andx  g02387(.a(n2466), .b(n2422), .O(n2552));
  andx  g02388(.a(n2424), .b(n2517), .O(n2553));
  orx   g02389(.a(n2553), .b(n2552), .O(n2554));
  andx  g02390(.a(n2554), .b(n2469), .O(n2555));
  orx   g02391(.a(n2424), .b(n2517), .O(n2556));
  orx   g02392(.a(n2466), .b(n2422), .O(n2557));
  andx  g02393(.a(n2557), .b(n2556), .O(n2558));
  andx  g02394(.a(n2558), .b(n2347), .O(n2559));
  orx   g02395(.a(n2559), .b(n2555), .O(n2560));
  andx  g02396(.a(n2515), .b(n2417), .O(n2561));
  andx  g02397(.a(n2420), .b(n2513), .O(n2562));
  orx   g02398(.a(n2562), .b(n2561), .O(n2563));
  andx  g02399(.a(n2563), .b(n2473), .O(n2564));
  orx   g02400(.a(n2420), .b(n2513), .O(n2565));
  orx   g02401(.a(n2515), .b(n2417), .O(n2566));
  andx  g02402(.a(n2566), .b(n2565), .O(n2567));
  andx  g02403(.a(n2567), .b(n2356), .O(n2568));
  orx   g02404(.a(n2568), .b(n2564), .O(n2569));
  orx   g02405(.a(n2414), .b(n2510), .O(n2570));
  orx   g02406(.a(n2475), .b(n2412), .O(n2571));
  andx  g02407(.a(n2571), .b(n2570), .O(n2572));
  orx   g02408(.a(n2572), .b(n2478), .O(n2573));
  andx  g02409(.a(n2475), .b(n2412), .O(n2574));
  andx  g02410(.a(n2414), .b(n2510), .O(n2575));
  orx   g02411(.a(n2575), .b(n2574), .O(n2576));
  orx   g02412(.a(n2576), .b(n2365), .O(n2577));
  andx  g02413(.a(n2577), .b(n2573), .O(n2578));
  andx  g02414(.a(n2400), .b(n2496), .O(n2579));
  orx   g02415(.a(n2579), .b(n2499), .O(n2580));
  orx   g02416(.a(n2501), .b(n2386), .O(n2581));
  orx   g02417(.a(n2581), .b(n2398), .O(n2582));
  andx  g02418(.a(n2582), .b(n2580), .O(n2583));
  orx   g02419(.a(n1766), .b(n1769), .O(n2584));
  andx  g02420(.a(n2584), .b(n1745), .O(n2585));
  orx   g02421(.a(n2585), .b(n2583), .O(n2586));
  orx   g02422(.a(n1793), .b(n254), .O(n2587));
  andx  g02423(.a(n2585), .b(n2583), .O(n2588));
  orx   g02424(.a(n2588), .b(n2587), .O(n2589));
  andx  g02425(.a(n2589), .b(n2586), .O(n2590));
  orx   g02426(.a(n2404), .b(n2503), .O(n2591));
  orx   g02427(.a(n2484), .b(n2402), .O(n2592));
  andx  g02428(.a(n2592), .b(n2591), .O(n2593));
  orx   g02429(.a(n2593), .b(n2377), .O(n2594));
  andx  g02430(.a(n2484), .b(n2402), .O(n2595));
  andx  g02431(.a(n2404), .b(n2503), .O(n2596));
  orx   g02432(.a(n2596), .b(n2595), .O(n2597));
  orx   g02433(.a(n2597), .b(n2487), .O(n2598));
  andx  g02434(.a(n2598), .b(n2594), .O(n2599));
  andx  g02435(.a(n2599), .b(n2590), .O(n2600));
  andx  g02436(.a(n1698), .b(n255), .O(n2601));
  invx  g02437(.a(n2601), .O(n2602));
  orx   g02438(.a(n2602), .b(n2600), .O(n2603));
  orx   g02439(.a(n2599), .b(n2590), .O(n2604));
  andx  g02440(.a(n2604), .b(n2603), .O(n2605));
  orx   g02441(.a(n2508), .b(n2407), .O(n2606));
  orx   g02442(.a(n2410), .b(n2506), .O(n2607));
  andx  g02443(.a(n2607), .b(n2606), .O(n2608));
  andx  g02444(.a(n2608), .b(n2482), .O(n2609));
  andx  g02445(.a(n2410), .b(n2506), .O(n2610));
  andx  g02446(.a(n2508), .b(n2407), .O(n2611));
  orx   g02447(.a(n2611), .b(n2610), .O(n2612));
  andx  g02448(.a(n2612), .b(n2372), .O(n2613));
  orx   g02449(.a(n2613), .b(n2609), .O(n2614));
  andx  g02450(.a(n2614), .b(n2605), .O(n2615));
  invx  g02451(.a(n2615), .O(n2616));
  andx  g02452(.a(n2581), .b(n2398), .O(n2617));
  andx  g02453(.a(n2579), .b(n2499), .O(n2618));
  orx   g02454(.a(n2618), .b(n2617), .O(n2619));
  andx  g02455(.a(n1774), .b(n1736), .O(n2620));
  orx   g02456(.a(n2620), .b(n1770), .O(n2621));
  andx  g02457(.a(n2621), .b(n2619), .O(n2622));
  andx  g02458(.a(n1559), .b(n255), .O(n2623));
  orx   g02459(.a(n2621), .b(n2619), .O(n2624));
  andx  g02460(.a(n2624), .b(n2623), .O(n2625));
  orx   g02461(.a(n2625), .b(n2622), .O(n2626));
  andx  g02462(.a(n2597), .b(n2487), .O(n2627));
  andx  g02463(.a(n2593), .b(n2377), .O(n2628));
  orx   g02464(.a(n2628), .b(n2627), .O(n2629));
  orx   g02465(.a(n2629), .b(n2626), .O(n2630));
  andx  g02466(.a(n2601), .b(n2630), .O(n2631));
  andx  g02467(.a(n2629), .b(n2626), .O(n2632));
  orx   g02468(.a(n2632), .b(n2631), .O(n2633));
  andx  g02469(.a(n1902), .b(n255), .O(n2634));
  orx   g02470(.a(n2634), .b(n2633), .O(n2635));
  orx   g02471(.a(n2612), .b(n2372), .O(n2636));
  orx   g02472(.a(n2608), .b(n2482), .O(n2637));
  andx  g02473(.a(n2637), .b(n2636), .O(n2638));
  orx   g02474(.a(n2634), .b(n2638), .O(n2639));
  andx  g02475(.a(n2639), .b(n2635), .O(n2640));
  andx  g02476(.a(n2640), .b(n2616), .O(n2641));
  andx  g02477(.a(n2641), .b(n2578), .O(n2642));
  orx   g02478(.a(n2641), .b(n2578), .O(n2643));
  andx  g02479(.a(n2116), .b(n255), .O(n2644));
  andx  g02480(.a(n2644), .b(n2643), .O(n2645));
  orx   g02481(.a(n2645), .b(n2642), .O(n2646));
  andx  g02482(.a(n2646), .b(n2569), .O(n2647));
  andx  g02483(.a(n2176), .b(n255), .O(n2648));
  orx   g02484(.a(n2646), .b(n2569), .O(n2649));
  andx  g02485(.a(n2649), .b(n2648), .O(n2650));
  orx   g02486(.a(n2650), .b(n2647), .O(n2651));
  orx   g02487(.a(n2558), .b(n2347), .O(n2654));
  orx   g02488(.a(n2554), .b(n2469), .O(n2655));
  andx  g02489(.a(n2655), .b(n2654), .O(n2656));
  invx  g02490(.a(n2647), .O(n2657));
  invx  g02491(.a(n2648), .O(n2658));
  orx   g02492(.a(n2567), .b(n2356), .O(n2659));
  orx   g02493(.a(n2563), .b(n2473), .O(n2660));
  andx  g02494(.a(n2660), .b(n2659), .O(n2661));
  invx  g02495(.a(n2642), .O(n2662));
  andx  g02496(.a(n2576), .b(n2365), .O(n2663));
  andx  g02497(.a(n2572), .b(n2478), .O(n2664));
  orx   g02498(.a(n2664), .b(n2663), .O(n2665));
  orx   g02499(.a(n1900), .b(n1823), .O(n2666));
  orx   g02500(.a(n1896), .b(n1824), .O(n2667));
  andx  g02501(.a(n2667), .b(n2666), .O(n2668));
  orx   g02502(.a(n2668), .b(n254), .O(n2669));
  andx  g02503(.a(n2669), .b(n2605), .O(n2670));
  andx  g02504(.a(n2669), .b(n2614), .O(n2671));
  orx   g02505(.a(n2671), .b(n2670), .O(n2672));
  orx   g02506(.a(n2672), .b(n2615), .O(n2673));
  andx  g02507(.a(n2673), .b(n2665), .O(n2674));
  invx  g02508(.a(n2644), .O(n2675));
  orx   g02509(.a(n2675), .b(n2674), .O(n2676));
  andx  g02510(.a(n2676), .b(n2662), .O(n2677));
  andx  g02511(.a(n2677), .b(n2661), .O(n2678));
  orx   g02512(.a(n2678), .b(n2658), .O(n2679));
  andx  g02513(.a(n2679), .b(n2657), .O(n2680));
  andx  g02514(.a(n2680), .b(n2656), .O(n2681));
  orx   g02515(.a(n254), .b(n2681), .O(n2684));
  orx   g02516(.a(n2651), .b(n2560), .O(n2687));
  andx  g02517(.a(n255), .b(n2687), .O(n2688));
  orx   g02518(.a(n2732), .b(n2532), .O(n2694));
  orx   g02519(.a(n2530), .b(n2527), .O(n2695));
  orx   g02520(.a(n2523), .b(n2338), .O(n2696));
  andx  g02521(.a(n2696), .b(n2695), .O(n2697));
  orx   g02522(.a(n2827), .b(n2697), .O(n2702));
  andx  g02523(.a(n2702), .b(n2694), .O(n2703));
  invx  g02524(.a(n1135), .O(n2704));
  andx  g02525(.a(n2535), .b(n2704), .O(n2705));
  andx  g02526(.a(n2429), .b(n2537), .O(n2722));
  orx   g02527(.a(n2722), .b(n2705), .O(n2723));
  invx  g02528(.a(n2723), .O(n2724));
  andx  g02529(.a(n255), .b(n2680), .O(n2730));
  andx  g02530(.a(n2730), .b(n2656), .O(n2732));
  orx   g02531(.a(n254), .b(n2651), .O(n2734));
  andx  g02532(.a(n2734), .b(n2560), .O(n2736));
  orx   g02533(.a(n2736), .b(n2732), .O(n2737));
  orx   g02534(.a(n2648), .b(n2677), .O(n2738));
  orx   g02535(.a(n2658), .b(n2646), .O(n2739));
  andx  g02536(.a(n2739), .b(n2738), .O(n2740));
  orx   g02537(.a(n2740), .b(n2661), .O(n2741));
  andx  g02538(.a(n2658), .b(n2646), .O(n2742));
  andx  g02539(.a(n2648), .b(n2677), .O(n2743));
  orx   g02540(.a(n2743), .b(n2742), .O(n2744));
  orx   g02541(.a(n2744), .b(n2569), .O(n2745));
  andx  g02542(.a(n2745), .b(n2741), .O(n2746));
  andx  g02543(.a(n2634), .b(n2633), .O(n2756));
  orx   g02544(.a(n2756), .b(n2670), .O(n2757));
  orx   g02545(.a(n2757), .b(n2614), .O(n2758));
  orx   g02546(.a(n2669), .b(n2605), .O(n2762));
  andx  g02547(.a(n2762), .b(n2635), .O(n2763));
  orx   g02548(.a(n2763), .b(n2638), .O(n2764));
  andx  g02549(.a(n2764), .b(n2758), .O(n2765));
  andx  g02550(.a(n2587), .b(n2621), .O(n2766));
  andx  g02551(.a(n2623), .b(n2585), .O(n2767));
  orx   g02552(.a(n2767), .b(n2766), .O(n2768));
  andx  g02553(.a(n2768), .b(n2583), .O(n2769));
  orx   g02554(.a(n2623), .b(n2585), .O(n2770));
  orx   g02555(.a(n2587), .b(n2621), .O(n2771));
  andx  g02556(.a(n2771), .b(n2770), .O(n2772));
  andx  g02557(.a(n2772), .b(n2619), .O(n2773));
  orx   g02558(.a(n2773), .b(n2769), .O(n2774));
  andx  g02559(.a(n1783), .b(n1718), .O(n2775));
  orx   g02560(.a(n1783), .b(n1718), .O(n2776));
  andx  g02561(.a(n2776), .b(n1714), .O(n2777));
  orx   g02562(.a(n2777), .b(n2775), .O(n2778));
  andx  g02563(.a(n2778), .b(n2774), .O(n2779));
  orx   g02564(.a(n2778), .b(n2774), .O(n2780));
  andx  g02565(.a(n1698), .b(n379), .O(n2781));
  andx  g02566(.a(n2781), .b(n2780), .O(n2782));
  orx   g02567(.a(n2782), .b(n2779), .O(n2783));
  andx  g02568(.a(n2783), .b(n1902), .O(n2784));
  andx  g02569(.a(n2602), .b(n2626), .O(n2785));
  andx  g02570(.a(n2601), .b(n2590), .O(n2786));
  orx   g02571(.a(n2786), .b(n2785), .O(n2787));
  andx  g02572(.a(n2787), .b(n2599), .O(n2788));
  orx   g02573(.a(n2601), .b(n2590), .O(n2789));
  orx   g02574(.a(n2602), .b(n2626), .O(n2790));
  andx  g02575(.a(n2790), .b(n2789), .O(n2791));
  andx  g02576(.a(n2791), .b(n2629), .O(n2792));
  orx   g02577(.a(n2792), .b(n2788), .O(n2793));
  andx  g02578(.a(n1902), .b(n379), .O(n2794));
  orx   g02579(.a(n2794), .b(n2783), .O(n2795));
  andx  g02580(.a(n2795), .b(n2793), .O(n2796));
  orx   g02581(.a(n2796), .b(n2784), .O(n2797));
  andx  g02582(.a(n2797), .b(n2765), .O(n2798));
  orx   g02583(.a(n2797), .b(n2765), .O(n2799));
  andx  g02584(.a(n2116), .b(n379), .O(n2800));
  andx  g02585(.a(n2800), .b(n2799), .O(n2801));
  orx   g02586(.a(n2801), .b(n2798), .O(n2802));
  andx  g02587(.a(n2802), .b(n2176), .O(n2803));
  andx  g02588(.a(n2644), .b(n2641), .O(n2804));
  andx  g02589(.a(n2675), .b(n2673), .O(n2805));
  orx   g02590(.a(n2805), .b(n2804), .O(n2806));
  orx   g02591(.a(n2806), .b(n2665), .O(n2807));
  orx   g02592(.a(n2675), .b(n2673), .O(n2808));
  orx   g02593(.a(n2644), .b(n2641), .O(n2809));
  andx  g02594(.a(n2809), .b(n2808), .O(n2810));
  orx   g02595(.a(n2810), .b(n2578), .O(n2811));
  andx  g02596(.a(n2811), .b(n2807), .O(n2812));
  andx  g02597(.a(n2176), .b(n379), .O(n2813));
  orx   g02598(.a(n2813), .b(n2802), .O(n2814));
  andx  g02599(.a(n2814), .b(n2812), .O(n2815));
  orx   g02600(.a(n2815), .b(n2803), .O(n2816));
  orx   g02601(.a(n2816), .b(n2746), .O(n2818));
  andx  g02602(.a(n379), .b(n2818), .O(n2821));
  orx   g02603(.a(n2734), .b(n2560), .O(n2827));
  orx   g02604(.a(n2730), .b(n2656), .O(n2828));
  andx  g02605(.a(n2828), .b(n2827), .O(n2829));
  andx  g02606(.a(n2744), .b(n2569), .O(n2831));
  andx  g02607(.a(n2740), .b(n2661), .O(n2832));
  orx   g02608(.a(n2832), .b(n2831), .O(n2833));
  andx  g02609(.a(n2763), .b(n2638), .O(n2834));
  andx  g02610(.a(n2757), .b(n2614), .O(n2835));
  orx   g02611(.a(n2835), .b(n2834), .O(n2836));
  orx   g02612(.a(n2772), .b(n2619), .O(n2837));
  orx   g02613(.a(n2768), .b(n2583), .O(n2838));
  andx  g02614(.a(n2838), .b(n2837), .O(n2839));
  orx   g02615(.a(n1776), .b(n1724), .O(n2840));
  andx  g02616(.a(n1776), .b(n1724), .O(n2841));
  orx   g02617(.a(n2841), .b(n1720), .O(n2842));
  andx  g02618(.a(n2842), .b(n2840), .O(n2843));
  orx   g02619(.a(n2843), .b(n2839), .O(n2844));
  andx  g02620(.a(n2843), .b(n2839), .O(n2845));
  orx   g02621(.a(n1696), .b(n1594), .O(n2846));
  orx   g02622(.a(n1692), .b(n1595), .O(n2847));
  andx  g02623(.a(n2847), .b(n2846), .O(n2848));
  orx   g02624(.a(n2848), .b(n378), .O(n2849));
  orx   g02625(.a(n2849), .b(n2845), .O(n2850));
  andx  g02626(.a(n2850), .b(n2844), .O(n2851));
  orx   g02627(.a(n2851), .b(n2668), .O(n2852));
  orx   g02628(.a(n2791), .b(n2629), .O(n2853));
  orx   g02629(.a(n2787), .b(n2599), .O(n2854));
  andx  g02630(.a(n2854), .b(n2853), .O(n2855));
  orx   g02631(.a(n2668), .b(n378), .O(n2856));
  andx  g02632(.a(n2856), .b(n2851), .O(n2857));
  orx   g02633(.a(n2857), .b(n2855), .O(n2858));
  andx  g02634(.a(n2858), .b(n2852), .O(n2859));
  orx   g02635(.a(n2859), .b(n2836), .O(n2860));
  andx  g02636(.a(n2859), .b(n2836), .O(n2861));
  orx   g02637(.a(n2114), .b(n2048), .O(n2862));
  orx   g02638(.a(n2107), .b(n2049), .O(n2863));
  andx  g02639(.a(n2863), .b(n2862), .O(n2864));
  orx   g02640(.a(n2864), .b(n378), .O(n2865));
  orx   g02641(.a(n2865), .b(n2861), .O(n2866));
  andx  g02642(.a(n2866), .b(n2860), .O(n2867));
  orx   g02643(.a(n2867), .b(n2333), .O(n2868));
  andx  g02644(.a(n2810), .b(n2578), .O(n2869));
  andx  g02645(.a(n2806), .b(n2665), .O(n2870));
  orx   g02646(.a(n2870), .b(n2869), .O(n2871));
  orx   g02647(.a(n2333), .b(n378), .O(n2872));
  andx  g02648(.a(n2872), .b(n2867), .O(n2873));
  orx   g02649(.a(n2873), .b(n2871), .O(n2874));
  andx  g02650(.a(n2874), .b(n2868), .O(n2875));
  andx  g02651(.a(n2875), .b(n2833), .O(n2876));
  orx   g02652(.a(n378), .b(n2876), .O(n2877));
  andx  g02653(.a(n2877), .b(n2829), .O(n2879));
  orx   g02654(.a(n2879), .b(n378), .O(n2880));
  orx   g02655(.a(n2821), .b(n2737), .O(n2883));
  andx  g02656(.a(n2883), .b(n379), .O(n2884));
  andx  g02657(.a(n2884), .b(n2703), .O(n2888));
  andx  g02658(.a(n2827), .b(n2697), .O(n2889));
  andx  g02659(.a(n2732), .b(n2532), .O(n2890));
  orx   g02660(.a(n2890), .b(n2889), .O(n2891));
  andx  g02661(.a(n2880), .b(n2891), .O(n2895));
  orx   g02662(.a(n2895), .b(n2888), .O(n2896));
  orx   g02663(.a(n378), .b(n2816), .O(n2899));
  andx  g02664(.a(n2899), .b(n2746), .O(n2900));
  andx  g02665(.a(n3185), .b(n2833), .O(n2904));
  orx   g02666(.a(n2904), .b(n2900), .O(n2905));
  andx  g02667(.a(n2176), .b(n250), .O(n2906));
  orx   g02668(.a(n2800), .b(n2797), .O(n2907));
  orx   g02669(.a(n2865), .b(n2859), .O(n2908));
  andx  g02670(.a(n2908), .b(n2907), .O(n2909));
  andx  g02671(.a(n2909), .b(n2836), .O(n2910));
  andx  g02672(.a(n2865), .b(n2859), .O(n2911));
  andx  g02673(.a(n2800), .b(n2797), .O(n2912));
  orx   g02674(.a(n2912), .b(n2911), .O(n2913));
  andx  g02675(.a(n2913), .b(n2765), .O(n2914));
  orx   g02676(.a(n2914), .b(n2910), .O(n2915));
  orx   g02677(.a(n2849), .b(n2843), .O(n2916));
  orx   g02678(.a(n2781), .b(n2778), .O(n2917));
  andx  g02679(.a(n2917), .b(n2916), .O(n2918));
  orx   g02680(.a(n2918), .b(n2774), .O(n2919));
  andx  g02681(.a(n2781), .b(n2778), .O(n2920));
  andx  g02682(.a(n2849), .b(n2843), .O(n2921));
  orx   g02683(.a(n2921), .b(n2920), .O(n2922));
  orx   g02684(.a(n2922), .b(n2839), .O(n2923));
  andx  g02685(.a(n2923), .b(n2919), .O(n2924));
  andx  g02686(.a(n1785), .b(n1699), .O(n2925));
  andx  g02687(.a(n1785), .b(n1593), .O(n2926));
  orx   g02688(.a(n2926), .b(n1700), .O(n2927));
  orx   g02689(.a(n2927), .b(n2925), .O(n2928));
  andx  g02690(.a(n2928), .b(n2924), .O(n2929));
  andx  g02691(.a(n1902), .b(n250), .O(n2930));
  andx  g02692(.a(n2930), .b(n2924), .O(n2931));
  andx  g02693(.a(n2930), .b(n2928), .O(n2932));
  orx   g02694(.a(n2932), .b(n2931), .O(n2933));
  orx   g02695(.a(n2933), .b(n2929), .O(n2934));
  andx  g02696(.a(n2116), .b(n250), .O(n2935));
  andx  g02697(.a(n2935), .b(n2934), .O(n2936));
  andx  g02698(.a(n2795), .b(n2852), .O(n2937));
  orx   g02699(.a(n2937), .b(n2793), .O(n2938));
  orx   g02700(.a(n2857), .b(n2784), .O(n2939));
  orx   g02701(.a(n2939), .b(n2855), .O(n2940));
  andx  g02702(.a(n2940), .b(n2938), .O(n2941));
  andx  g02703(.a(n2941), .b(n2934), .O(n2942));
  andx  g02704(.a(n2941), .b(n2935), .O(n2943));
  orx   g02705(.a(n2943), .b(n2942), .O(n2944));
  orx   g02706(.a(n2944), .b(n2936), .O(n2945));
  andx  g02707(.a(n2945), .b(n2915), .O(n2946));
  orx   g02708(.a(n2946), .b(n2906), .O(n2947));
  orx   g02709(.a(n2913), .b(n2765), .O(n2948));
  orx   g02710(.a(n2909), .b(n2836), .O(n2949));
  andx  g02711(.a(n2949), .b(n2948), .O(n2950));
  andx  g02712(.a(n2922), .b(n2839), .O(n2951));
  andx  g02713(.a(n2918), .b(n2774), .O(n2952));
  orx   g02714(.a(n2952), .b(n2951), .O(n2953));
  andx  g02715(.a(n1783), .b(n1780), .O(n2954));
  andx  g02716(.a(n1776), .b(n1726), .O(n2955));
  orx   g02717(.a(n2955), .b(n2954), .O(n2956));
  orx   g02718(.a(n2956), .b(n1711), .O(n2957));
  orx   g02719(.a(n1711), .b(n1710), .O(n2958));
  orx   g02720(.a(n2956), .b(n1710), .O(n2959));
  andx  g02721(.a(n2959), .b(n2958), .O(n2960));
  andx  g02722(.a(n2960), .b(n2957), .O(n2961));
  orx   g02723(.a(n2961), .b(n2953), .O(n2962));
  invx  g02724(.a(n2930), .O(n2963));
  orx   g02725(.a(n2963), .b(n2953), .O(n2964));
  orx   g02726(.a(n2963), .b(n2961), .O(n2965));
  andx  g02727(.a(n2965), .b(n2964), .O(n2966));
  andx  g02728(.a(n2966), .b(n2962), .O(n2967));
  orx   g02729(.a(n2864), .b(n179), .O(n2968));
  orx   g02730(.a(n2968), .b(n2967), .O(n2969));
  andx  g02731(.a(n2939), .b(n2855), .O(n2970));
  andx  g02732(.a(n2937), .b(n2793), .O(n2971));
  orx   g02733(.a(n2971), .b(n2970), .O(n2972));
  orx   g02734(.a(n2972), .b(n2967), .O(n2973));
  orx   g02735(.a(n2972), .b(n2968), .O(n2974));
  andx  g02736(.a(n2974), .b(n2973), .O(n2975));
  andx  g02737(.a(n2975), .b(n2969), .O(n2976));
  andx  g02738(.a(n2976), .b(n2950), .O(n2977));
  invx  g02739(.a(n2977), .O(n2978));
  andx  g02740(.a(n2978), .b(n2947), .O(n2979));
  orx   g02741(.a(n2873), .b(n2803), .O(n2980));
  andx  g02742(.a(n2980), .b(n2812), .O(n2981));
  andx  g02743(.a(n2814), .b(n2868), .O(n2982));
  andx  g02744(.a(n2982), .b(n2871), .O(n2983));
  orx   g02745(.a(n2983), .b(n2981), .O(n2984));
  andx  g02746(.a(n250), .b(n2984), .O(n2989));
  orx   g02747(.a(n2989), .b(n2979), .O(n2990));
  andx  g02748(.a(n250), .b(n2905), .O(n2994));
  orx   g02749(.a(n2990), .b(n2994), .O(n2996));
  andx  g02750(.a(n2904), .b(n2829), .O(n3001));
  andx  g02751(.a(n3014), .b(n2737), .O(n3005));
  orx   g02752(.a(n3005), .b(n3001), .O(n3006));
  andx  g02753(.a(n3006), .b(n2996), .O(n3007));
  invx  g02754(.a(n3007), .O(n3008));
  orx   g02755(.a(n2723), .b(n179), .O(n3011));
  orx   g02756(.a(n3185), .b(n2833), .O(n3013));
  orx   g02757(.a(n2899), .b(n2746), .O(n3014));
  andx  g02758(.a(n3014), .b(n3013), .O(n3015));
  orx   g02759(.a(n179), .b(n3015), .O(n3017));
  orx   g02760(.a(n2333), .b(n179), .O(n3018));
  orx   g02761(.a(n2976), .b(n2950), .O(n3019));
  andx  g02762(.a(n3019), .b(n3018), .O(n3020));
  orx   g02763(.a(n2977), .b(n3020), .O(n3021));
  orx   g02764(.a(n2982), .b(n2871), .O(n3022));
  orx   g02765(.a(n2980), .b(n2812), .O(n3023));
  andx  g02766(.a(n3023), .b(n3022), .O(n3024));
  orx   g02767(.a(n179), .b(n3024), .O(n3027));
  andx  g02768(.a(n3027), .b(n3021), .O(n3028));
  andx  g02769(.a(n3028), .b(n3017), .O(n3031));
  orx   g02770(.a(n3014), .b(n2737), .O(n3033));
  orx   g02771(.a(n2904), .b(n2829), .O(n3034));
  andx  g02772(.a(n3034), .b(n3033), .O(n3035));
  orx   g02773(.a(n3008), .b(n2896), .O(n3039));
  andx  g02774(.a(n2176), .b(n554), .O(n3040));
  invx  g02775(.a(n3040), .O(n3041));
  andx  g02776(.a(n2121), .b(n1967), .O(n3042));
  invx  g02777(.a(n3042), .O(n3043));
  andx  g02778(.a(n2047), .b(n2127), .O(n3044));
  orx   g02779(.a(n3044), .b(n2122), .O(n3045));
  andx  g02780(.a(n3045), .b(n3043), .O(n3046));
  orx   g02781(.a(n3046), .b(n3041), .O(n3047));
  orx   g02782(.a(n2121), .b(n1967), .O(n3048));
  andx  g02783(.a(n3048), .b(n2117), .O(n3049));
  orx   g02784(.a(n3049), .b(n3042), .O(n3050));
  orx   g02785(.a(n3050), .b(n3040), .O(n3051));
  andx  g02786(.a(n3051), .b(n3047), .O(n3052));
  andx  g02787(.a(n1816), .b(n1559), .O(n3053));
  invx  g02788(.a(n3053), .O(n3054));
  andx  g02789(.a(n1812), .b(n1793), .O(n3055));
  orx   g02790(.a(n3055), .b(n1814), .O(n3056));
  andx  g02791(.a(n3056), .b(n3054), .O(n3057));
  andx  g02792(.a(n1902), .b(n836), .O(n3058));
  invx  g02793(.a(n3058), .O(n3059));
  andx  g02794(.a(n3059), .b(n3057), .O(n3060));
  invx  g02795(.a(n3057), .O(n3061));
  andx  g02796(.a(n3058), .b(n3061), .O(n3062));
  orx   g02797(.a(n3062), .b(n3060), .O(n3063));
  invx  g02798(.a(n3063), .O(n3064));
  andx  g02799(.a(n3064), .b(n2848), .O(n3065));
  andx  g02800(.a(n3063), .b(n1698), .O(n3066));
  orx   g02801(.a(n3066), .b(n3065), .O(n3067));
  andx  g02802(.a(n1959), .b(n1822), .O(n3068));
  orx   g02803(.a(n1959), .b(n1822), .O(n3069));
  andx  g02804(.a(n3069), .b(n1903), .O(n3070));
  orx   g02805(.a(n3070), .b(n3068), .O(n3071));
  andx  g02806(.a(n3071), .b(n2116), .O(n3072));
  invx  g02807(.a(n3072), .O(n3073));
  andx  g02808(.a(n2116), .b(n605), .O(n3074));
  orx   g02809(.a(n3074), .b(n3071), .O(n3075));
  andx  g02810(.a(n3075), .b(n3073), .O(n3076));
  orx   g02811(.a(n3076), .b(n3067), .O(n3077));
  andx  g02812(.a(n3076), .b(n3067), .O(n3078));
  invx  g02813(.a(n3078), .O(n3079));
  andx  g02814(.a(n3079), .b(n3077), .O(n3080));
  andx  g02815(.a(n3080), .b(n3052), .O(n3081));
  andx  g02816(.a(n3050), .b(n3040), .O(n3082));
  andx  g02817(.a(n3046), .b(n3041), .O(n3083));
  orx   g02818(.a(n3083), .b(n3082), .O(n3084));
  invx  g02819(.a(n3080), .O(n3085));
  andx  g02820(.a(n3085), .b(n3084), .O(n3086));
  orx   g02821(.a(n3086), .b(n3081), .O(n3087));
  andx  g02822(.a(n2335), .b(n2330), .O(n3088));
  orx   g02823(.a(n3088), .b(n2293), .O(n3089));
  orx   g02824(.a(n2325), .b(n2132), .O(n3091));
  andx  g02825(.a(n3091), .b(n2334), .O(n3092));
  orx   g02826(.a(n477), .b(n3089), .O(n3096));
  andx  g02827(.a(n3096), .b(n3087), .O(n3097));
  orx   g02828(.a(n3085), .b(n3084), .O(n3098));
  orx   g02829(.a(n3080), .b(n3052), .O(n3099));
  andx  g02830(.a(n3099), .b(n3098), .O(n3100));
  andx  g02831(.a(n488), .b(n3092), .O(n3103));
  andx  g02832(.a(n3103), .b(n3100), .O(n3104));
  orx   g02833(.a(n3104), .b(n3097), .O(n3105));
  orx   g02834(.a(n2427), .b(n2527), .O(n3107));
  andx  g02835(.a(n3107), .b(n499), .O(n3108));
  andx  g02836(.a(n2520), .b(n2338), .O(n3113));
  orx   g02837(.a(n3113), .b(n481), .O(n3114));
  andx  g02838(.a(n2524), .b(n3105), .O(n3119));
  orx   g02839(.a(n3103), .b(n3100), .O(n3120));
  orx   g02840(.a(n3096), .b(n3087), .O(n3121));
  andx  g02841(.a(n3121), .b(n3120), .O(n3122));
  andx  g02842(.a(n2695), .b(n3122), .O(n3126));
  orx   g02843(.a(n3126), .b(n3119), .O(n3127));
  orx   g02844(.a(n254), .b(n2697), .O(n3128));
  andx  g02845(.a(n3128), .b(n2684), .O(n3129));
  andx  g02846(.a(n255), .b(n2532), .O(n3131));
  orx   g02847(.a(n3131), .b(n2688), .O(n3132));
  orx   g02848(.a(n3132), .b(n3127), .O(n3136));
  orx   g02849(.a(n2695), .b(n3122), .O(n3137));
  orx   g02850(.a(n2524), .b(n3105), .O(n3138));
  andx  g02851(.a(n3138), .b(n3137), .O(n3139));
  orx   g02852(.a(n3129), .b(n3139), .O(n3144));
  andx  g02853(.a(n3144), .b(n3136), .O(n3145));
  orx   g02854(.a(n3159), .b(n3145), .O(n3151));
  andx  g02855(.a(n3129), .b(n3139), .O(n3152));
  andx  g02856(.a(n3132), .b(n3127), .O(n3153));
  orx   g02857(.a(n3153), .b(n3152), .O(n3154));
  orx   g02858(.a(n2888), .b(n3154), .O(n3156));
  andx  g02859(.a(n3156), .b(n3151), .O(n3157));
  orx   g02860(.a(n3157), .b(n3039), .O(n3158));
  orx   g02861(.a(n2880), .b(n2891), .O(n3159));
  orx   g02862(.a(n2884), .b(n2703), .O(n3160));
  andx  g02863(.a(n3160), .b(n3159), .O(n3161));
  andx  g02864(.a(n3007), .b(n3161), .O(n3166));
  andx  g02865(.a(n2888), .b(n3154), .O(n3167));
  andx  g02866(.a(n3159), .b(n3145), .O(n3168));
  orx   g02867(.a(n3168), .b(n3167), .O(n3169));
  orx   g02868(.a(n3169), .b(n3166), .O(n3170));
  andx  g02869(.a(n3170), .b(n3158), .O(n3171));
  andx  g02870(.a(n3031), .b(n3006), .O(n3175));
  andx  g02871(.a(n2996), .b(n3035), .O(n3179));
  orx   g02872(.a(n3179), .b(n3175), .O(n3180));
  orx   g02873(.a(n2996), .b(n3035), .O(n3181));
  orx   g02874(.a(n3031), .b(n3006), .O(n3182));
  andx  g02875(.a(n3182), .b(n3181), .O(n3183));
  andx  g02876(.a(n379), .b(n2875), .O(n3185));
  andx  g02877(.a(n3269), .b(n3015), .O(n3194));
  andx  g02878(.a(n3209), .b(n2905), .O(n3200));
  orx   g02879(.a(n3200), .b(n3194), .O(n3201));
  orx   g02880(.a(n179), .b(n2979), .O(n3202));
  andx  g02881(.a(n3202), .b(n2984), .O(n3205));
  andx  g02882(.a(n250), .b(n3021), .O(n3206));
  andx  g02883(.a(n3206), .b(n3024), .O(n3209));
  orx   g02884(.a(n3209), .b(n3205), .O(n3210));
  andx  g02885(.a(n3210), .b(n827), .O(n3211));
  invx  g02886(.a(n3211), .O(n3212));
  andx  g02887(.a(n2976), .b(n3018), .O(n3213));
  andx  g02888(.a(n2945), .b(n2906), .O(n3214));
  orx   g02889(.a(n3214), .b(n3213), .O(n3215));
  andx  g02890(.a(n3215), .b(n2915), .O(n3216));
  orx   g02891(.a(n2945), .b(n2906), .O(n3217));
  orx   g02892(.a(n2976), .b(n3018), .O(n3218));
  andx  g02893(.a(n3218), .b(n3217), .O(n3219));
  andx  g02894(.a(n3219), .b(n2950), .O(n3220));
  orx   g02895(.a(n3220), .b(n3216), .O(n3221));
  orx   g02896(.a(n2968), .b(n2934), .O(n3222));
  orx   g02897(.a(n2935), .b(n2967), .O(n3223));
  andx  g02898(.a(n3223), .b(n3222), .O(n3224));
  andx  g02899(.a(n3224), .b(n2941), .O(n3225));
  andx  g02900(.a(n2935), .b(n2967), .O(n3226));
  andx  g02901(.a(n2968), .b(n2934), .O(n3227));
  orx   g02902(.a(n3227), .b(n3226), .O(n3228));
  andx  g02903(.a(n3228), .b(n2972), .O(n3229));
  orx   g02904(.a(n3229), .b(n3225), .O(n3230));
  andx  g02905(.a(n3230), .b(n827), .O(n3231));
  andx  g02906(.a(n3231), .b(n3221), .O(n3232));
  invx  g02907(.a(n3232), .O(n3233));
  orx   g02908(.a(n3219), .b(n2950), .O(n3234));
  orx   g02909(.a(n3215), .b(n2915), .O(n3235));
  andx  g02910(.a(n3235), .b(n3234), .O(n3236));
  orx   g02911(.a(n3228), .b(n2972), .O(n3237));
  orx   g02912(.a(n3224), .b(n2941), .O(n3238));
  andx  g02913(.a(n3238), .b(n3237), .O(n3239));
  andx  g02914(.a(n3239), .b(n3236), .O(n3240));
  andx  g02915(.a(n1790), .b(n827), .O(n3241));
  andx  g02916(.a(n2963), .b(n2928), .O(n3242));
  andx  g02917(.a(n2930), .b(n2961), .O(n3243));
  orx   g02918(.a(n3243), .b(n3242), .O(n3244));
  orx   g02919(.a(n2924), .b(n3244), .O(n3253));
  orx   g02920(.a(n2930), .b(n2961), .O(n3254));
  orx   g02921(.a(n2963), .b(n2928), .O(n3255));
  andx  g02922(.a(n3255), .b(n3254), .O(n3256));
  orx   g02923(.a(n2953), .b(n3256), .O(n3257));
  andx  g02924(.a(n3257), .b(n3253), .O(n3258));
  andx  g02925(.a(n3258), .b(n3241), .O(n3259));
  andx  g02926(.a(n3258), .b(n3231), .O(n3260));
  orx   g02927(.a(n3260), .b(n3259), .O(n3261));
  invx  g02928(.a(n3261), .O(n3262));
  orx   g02929(.a(n3262), .b(n3240), .O(n3263));
  andx  g02930(.a(n3263), .b(n3233), .O(n3264));
  invx  g02931(.a(n3264), .O(n3265));
  andx  g02932(.a(n3265), .b(n3221), .O(n3266));
  invx  g02933(.a(n3266), .O(n3267));
  orx   g02934(.a(n3206), .b(n3024), .O(n3268));
  orx   g02935(.a(n3202), .b(n2984), .O(n3269));
  andx  g02936(.a(n3269), .b(n3268), .O(n3270));
  andx  g02937(.a(n3221), .b(n827), .O(n3271));
  invx  g02938(.a(n3271), .O(n3272));
  andx  g02939(.a(n3272), .b(n3264), .O(n3273));
  orx   g02940(.a(n3273), .b(n3270), .O(n3274));
  andx  g02941(.a(n3274), .b(n3267), .O(n3275));
  andx  g02942(.a(n3275), .b(n3212), .O(n3276));
  orx   g02943(.a(n3276), .b(n3201), .O(n3277));
  invx  g02944(.a(n3275), .O(n3278));
  andx  g02945(.a(n3274), .b(n3277), .O(n3281));
  orx   g02946(.a(n3209), .b(n2905), .O(n3282));
  orx   g02947(.a(n3269), .b(n3015), .O(n3283));
  andx  g02948(.a(n3283), .b(n3282), .O(n3284));
  andx  g02949(.a(n3284), .b(n827), .O(n3285));
  invx  g02950(.a(n3285), .O(n3286));
  andx  g02951(.a(n3286), .b(n3281), .O(n3287));
  orx   g02952(.a(n3287), .b(n3183), .O(n3288));
  invx  g02953(.a(n3281), .O(n3289));
  andx  g02954(.a(n3277), .b(n3288), .O(n3292));
  invx  g02955(.a(n3292), .O(n3293));
  andx  g02956(.a(n3008), .b(n2896), .O(n3296));
  orx   g02957(.a(n3296), .b(n3166), .O(n3297));
  andx  g02958(.a(n3180), .b(n827), .O(n3298));
  invx  g02959(.a(n3298), .O(n3299));
  andx  g02960(.a(n3299), .b(n3292), .O(n3300));
  orx   g02961(.a(n3300), .b(n3297), .O(n3301));
  andx  g02962(.a(n3301), .b(n3288), .O(n3302));
  invx  g02963(.a(n3302), .O(n3303));
  andx  g02964(.a(n3303), .b(n3171), .O(n3304));
  invx  g02965(.a(n3304), .O(n3305));
  andx  g02966(.a(n3171), .b(n827), .O(n3306));
  invx  g02967(.a(n3306), .O(n3307));
  andx  g02968(.a(n3307), .b(n3302), .O(n3308));
  orx   g02969(.a(n3308), .b(n3297), .O(n3309));
  andx  g02970(.a(n3309), .b(n3305), .O(n3310));
  invx  g02971(.a(n3310), .O(n3311));
  andx  g02972(.a(n2888), .b(n3145), .O(n3312));
  invx  g02973(.a(n3312), .O(n3313));
  andx  g02974(.a(n3057), .b(n2848), .O(n3318));
  orx   g02975(.a(n3318), .b(n3059), .O(n3319));
  andx  g02976(.a(n3319), .b(n3056), .O(n3320));
  andx  g02977(.a(n2116), .b(n836), .O(n3321));
  invx  g02978(.a(n3321), .O(n3322));
  andx  g02979(.a(n3322), .b(n3320), .O(n3323));
  invx  g02980(.a(n3320), .O(n3324));
  andx  g02981(.a(n3321), .b(n3324), .O(n3325));
  orx   g02982(.a(n3325), .b(n3323), .O(n3326));
  invx  g02983(.a(n3326), .O(n3327));
  andx  g02984(.a(n3327), .b(n2668), .O(n3328));
  andx  g02985(.a(n3326), .b(n1902), .O(n3329));
  orx   g02986(.a(n3329), .b(n3328), .O(n3330));
  invx  g02987(.a(n3330), .O(n3331));
  andx  g02988(.a(n3075), .b(n3067), .O(n3332));
  orx   g02989(.a(n3332), .b(n3072), .O(n3333));
  andx  g02990(.a(n3333), .b(n2176), .O(n3334));
  invx  g02991(.a(n3334), .O(n3335));
  andx  g02992(.a(n2176), .b(n605), .O(n3336));
  orx   g02993(.a(n3336), .b(n3333), .O(n3337));
  andx  g02994(.a(n3337), .b(n3335), .O(n3338));
  invx  g02995(.a(n3338), .O(n3339));
  andx  g02996(.a(n3339), .b(n3331), .O(n3340));
  andx  g02997(.a(n3338), .b(n3330), .O(n3341));
  orx   g02998(.a(n3341), .b(n3340), .O(n3342));
  andx  g02999(.a(n3080), .b(n3050), .O(n3345));
  invx  g03000(.a(n3345), .O(n3346));
  andx  g03001(.a(n3085), .b(n3046), .O(n3347));
  orx   g03002(.a(n3347), .b(n3041), .O(n3348));
  andx  g03003(.a(n3348), .b(n3346), .O(n3349));
  andx  g03004(.a(n554), .b(n3349), .O(n3353));
  andx  g03005(.a(n3353), .b(n3342), .O(n3354));
  invx  g03006(.a(n3342), .O(n3355));
  orx   g03007(.a(n560), .b(n3593), .O(n3357));
  andx  g03008(.a(n3357), .b(n3355), .O(n3358));
  orx   g03009(.a(n3358), .b(n3354), .O(n3359));
  andx  g03010(.a(n488), .b(n3100), .O(n3360));
  orx   g03011(.a(n3360), .b(n3089), .O(n3361));
  invx  g03012(.a(n3361), .O(n3363));
  andx  g03013(.a(n488), .b(n3363), .O(n3366));
  orx   g03014(.a(n3366), .b(n3359), .O(n3367));
  orx   g03015(.a(n3357), .b(n3355), .O(n3368));
  orx   g03016(.a(n3353), .b(n3342), .O(n3369));
  andx  g03017(.a(n3369), .b(n3368), .O(n3370));
  orx   g03018(.a(n477), .b(n3361), .O(n3372));
  orx   g03019(.a(n3372), .b(n3370), .O(n3373));
  andx  g03020(.a(n3373), .b(n3367), .O(n3374));
  andx  g03021(.a(n3114), .b(n3105), .O(n3379));
  orx   g03022(.a(n3379), .b(n481), .O(n3380));
  orx   g03023(.a(n3108), .b(n3122), .O(n3383));
  andx  g03024(.a(n3383), .b(n499), .O(n3384));
  andx  g03025(.a(n3384), .b(n3374), .O(n3388));
  andx  g03026(.a(n3372), .b(n3370), .O(n3389));
  andx  g03027(.a(n3366), .b(n3359), .O(n3390));
  orx   g03028(.a(n3390), .b(n3389), .O(n3391));
  andx  g03029(.a(n3380), .b(n3391), .O(n3395));
  orx   g03030(.a(n3395), .b(n3388), .O(n3396));
  orx   g03031(.a(n3396), .b(n3153), .O(n3397));
  orx   g03032(.a(n3380), .b(n3391), .O(n3399));
  orx   g03033(.a(n3384), .b(n3374), .O(n3400));
  andx  g03034(.a(n3400), .b(n3399), .O(n3401));
  orx   g03035(.a(n3401), .b(n3144), .O(n3402));
  andx  g03036(.a(n3402), .b(n3397), .O(n3403));
  orx   g03037(.a(n3403), .b(n3313), .O(n3404));
  orx   g03038(.a(n3403), .b(n3158), .O(n3405));
  andx  g03039(.a(n3405), .b(n3404), .O(n3406));
  andx  g03040(.a(n3169), .b(n3166), .O(n3407));
  andx  g03041(.a(n3401), .b(n3144), .O(n3408));
  andx  g03042(.a(n3396), .b(n3153), .O(n3409));
  orx   g03043(.a(n3409), .b(n3408), .O(n3410));
  orx   g03044(.a(n3410), .b(n3312), .O(n3411));
  orx   g03045(.a(n3411), .b(n3407), .O(n3412));
  andx  g03046(.a(n3412), .b(n3406), .O(n3413));
  andx  g03047(.a(n3413), .b(n827), .O(n3414));
  invx  g03048(.a(n3414), .O(n3415));
  andx  g03049(.a(n3415), .b(n3171), .O(n3416));
  andx  g03050(.a(n3157), .b(n3039), .O(n3417));
  orx   g03051(.a(n3417), .b(n3407), .O(n3418));
  andx  g03052(.a(n3414), .b(n3418), .O(n3419));
  orx   g03053(.a(n3419), .b(n3416), .O(n3420));
  andx  g03054(.a(n3420), .b(n3311), .O(n3421));
  invx  g03055(.a(n3421), .O(n3422));
  orx   g03056(.a(n3420), .b(n3311), .O(n3423));
  andx  g03057(.a(n3423), .b(n3422), .O(n3424));
  invx  g03058(.a(n3424), .O(n3425));
  andx  g03059(.a(n3297), .b(n827), .O(n3426));
  andx  g03060(.a(n3426), .b(n3171), .O(n3427));
  orx   g03061(.a(n3007), .b(n3161), .O(n3428));
  andx  g03062(.a(n3428), .b(n3039), .O(n3429));
  andx  g03063(.a(n3307), .b(n3429), .O(n3430));
  orx   g03064(.a(n3430), .b(n3427), .O(n3431));
  andx  g03065(.a(n3431), .b(n3303), .O(n3432));
  invx  g03066(.a(n3432), .O(n3433));
  orx   g03067(.a(n3431), .b(n3303), .O(n3434));
  andx  g03068(.a(n3434), .b(n3433), .O(n3435));
  andx  g03069(.a(n3429), .b(n827), .O(n3436));
  orx   g03070(.a(n3436), .b(n3183), .O(n3437));
  andx  g03071(.a(n3183), .b(n827), .O(n3438));
  andx  g03072(.a(n3438), .b(n3429), .O(n3439));
  invx  g03073(.a(n3439), .O(n3440));
  andx  g03074(.a(n3440), .b(n3437), .O(n3441));
  invx  g03075(.a(n3441), .O(n3442));
  andx  g03076(.a(n3442), .b(n3293), .O(n3443));
  andx  g03077(.a(n3441), .b(n3292), .O(n3444));
  orx   g03078(.a(n3444), .b(n3443), .O(n3445));
  invx  g03079(.a(n3445), .O(n3446));
  andx  g03080(.a(n3299), .b(n3284), .O(n3447));
  andx  g03081(.a(n3201), .b(n827), .O(n3448));
  andx  g03082(.a(n3448), .b(n3180), .O(n3449));
  orx   g03083(.a(n3449), .b(n3447), .O(n3450));
  andx  g03084(.a(n3450), .b(n3289), .O(n3451));
  invx  g03085(.a(n3451), .O(n3452));
  orx   g03086(.a(n3450), .b(n3289), .O(n3453));
  andx  g03087(.a(n3453), .b(n3452), .O(n3454));
  andx  g03088(.a(n3270), .b(n827), .O(n3455));
  andx  g03089(.a(n3455), .b(n3284), .O(n3456));
  andx  g03090(.a(n3286), .b(n3210), .O(n3457));
  orx   g03091(.a(n3457), .b(n3456), .O(n3458));
  andx  g03092(.a(n3458), .b(n3278), .O(n3459));
  invx  g03093(.a(n3459), .O(n3460));
  orx   g03094(.a(n3458), .b(n3278), .O(n3461));
  andx  g03095(.a(n3461), .b(n3460), .O(n3462));
  andx  g03096(.a(n3236), .b(n3211), .O(n3463));
  andx  g03097(.a(n3221), .b(n3270), .O(n3464));
  andx  g03098(.a(n3221), .b(n826), .O(n3465));
  orx   g03099(.a(n3465), .b(n3464), .O(n3466));
  orx   g03100(.a(n3466), .b(n3463), .O(n3467));
  andx  g03101(.a(n3467), .b(n3264), .O(n3468));
  invx  g03102(.a(n3468), .O(n3469));
  orx   g03103(.a(n3467), .b(n3264), .O(n3470));
  andx  g03104(.a(n3470), .b(n3469), .O(n3471));
  invx  g03105(.a(n3471), .O(n3472));
  andx  g03106(.a(n3210), .b(n299), .O(n3473));
  andx  g03107(.a(n3258), .b(n299), .O(n3474));
  andx  g03108(.a(n3474), .b(n3241), .O(n3475));
  andx  g03109(.a(n3230), .b(n299), .O(n3476));
  andx  g03110(.a(n3476), .b(n3475), .O(n3477));
  andx  g03111(.a(n1789), .b(n827), .O(n3478));
  andx  g03112(.a(n3478), .b(n3258), .O(n3479));
  invx  g03113(.a(n3479), .O(n3480));
  andx  g03114(.a(n3258), .b(n827), .O(n3481));
  orx   g03115(.a(n3481), .b(n1789), .O(n3482));
  andx  g03116(.a(n3482), .b(n3480), .O(n3483));
  invx  g03117(.a(n3483), .O(n3484));
  andx  g03118(.a(n3484), .b(n3476), .O(n3485));
  orx   g03119(.a(n3485), .b(n3477), .O(n3486));
  andx  g03120(.a(n3486), .b(n3221), .O(n3487));
  andx  g03121(.a(n2953), .b(n3256), .O(n3488));
  andx  g03122(.a(n2924), .b(n3244), .O(n3489));
  orx   g03123(.a(n3489), .b(n3488), .O(n3490));
  invx  g03124(.a(n3231), .O(n3491));
  invx  g03125(.a(n3259), .O(n3492));
  andx  g03126(.a(n3492), .b(n3491), .O(n3493));
  andx  g03127(.a(n3259), .b(n3231), .O(n3494));
  orx   g03128(.a(n3494), .b(n3493), .O(n3495));
  andx  g03129(.a(n3495), .b(n3490), .O(n3496));
  invx  g03130(.a(n3496), .O(n3497));
  orx   g03131(.a(n3495), .b(n3490), .O(n3498));
  andx  g03132(.a(n3498), .b(n3497), .O(n3499));
  andx  g03133(.a(n3221), .b(n299), .O(n3500));
  orx   g03134(.a(n3500), .b(n3486), .O(n3501));
  andx  g03135(.a(n3501), .b(n3499), .O(n3502));
  orx   g03136(.a(n3502), .b(n3487), .O(n3503));
  andx  g03137(.a(n3503), .b(n3473), .O(n3504));
  invx  g03138(.a(n3504), .O(n3505));
  andx  g03139(.a(n3272), .b(n3239), .O(n3506));
  orx   g03140(.a(n3506), .b(n3232), .O(n3507));
  andx  g03141(.a(n3507), .b(n3261), .O(n3508));
  invx  g03142(.a(n3508), .O(n3509));
  orx   g03143(.a(n3507), .b(n3261), .O(n3510));
  andx  g03144(.a(n3510), .b(n3509), .O(n3511));
  invx  g03145(.a(n3473), .O(n3512));
  invx  g03146(.a(n3503), .O(n3513));
  andx  g03147(.a(n3513), .b(n3512), .O(n3514));
  orx   g03148(.a(n3514), .b(n3511), .O(n3515));
  andx  g03149(.a(n3515), .b(n3505), .O(n3516));
  invx  g03150(.a(n3516), .O(n3517));
  andx  g03151(.a(n3517), .b(n3472), .O(n3518));
  invx  g03152(.a(n3518), .O(n3519));
  andx  g03153(.a(n3516), .b(n3471), .O(n3520));
  andx  g03154(.a(n3284), .b(n299), .O(n3521));
  invx  g03155(.a(n3521), .O(n3522));
  orx   g03156(.a(n3522), .b(n3520), .O(n3523));
  andx  g03157(.a(n3523), .b(n3519), .O(n3524));
  invx  g03158(.a(n3524), .O(n3525));
  andx  g03159(.a(n3525), .b(n3462), .O(n3526));
  invx  g03160(.a(n3526), .O(n3527));
  andx  g03161(.a(n3180), .b(n299), .O(n3528));
  invx  g03162(.a(n3528), .O(n3529));
  invx  g03163(.a(n3462), .O(n3530));
  andx  g03164(.a(n3524), .b(n3530), .O(n3531));
  orx   g03165(.a(n3531), .b(n3529), .O(n3532));
  andx  g03166(.a(n3532), .b(n3527), .O(n3533));
  invx  g03167(.a(n3533), .O(n3534));
  andx  g03168(.a(n3534), .b(n3454), .O(n3535));
  invx  g03169(.a(n3535), .O(n3536));
  andx  g03170(.a(n3429), .b(n299), .O(n3537));
  invx  g03171(.a(n3537), .O(n3538));
  invx  g03172(.a(n3454), .O(n3539));
  andx  g03173(.a(n3533), .b(n3539), .O(n3540));
  orx   g03174(.a(n3540), .b(n3538), .O(n3541));
  andx  g03175(.a(n3541), .b(n3536), .O(n3542));
  invx  g03176(.a(n3542), .O(n3543));
  andx  g03177(.a(n3543), .b(n3446), .O(n3544));
  invx  g03178(.a(n3544), .O(n3545));
  andx  g03179(.a(n3171), .b(n299), .O(n3546));
  invx  g03180(.a(n3546), .O(n3547));
  andx  g03181(.a(n3542), .b(n3445), .O(n3548));
  orx   g03182(.a(n3548), .b(n3547), .O(n3549));
  andx  g03183(.a(n3549), .b(n3545), .O(n3550));
  invx  g03184(.a(n3550), .O(n3551));
  andx  g03185(.a(n3551), .b(n3435), .O(n3552));
  invx  g03186(.a(n3552), .O(n3553));
  andx  g03187(.a(n3413), .b(n299), .O(n3554));
  invx  g03188(.a(n3554), .O(n3555));
  invx  g03189(.a(n3435), .O(n3556));
  andx  g03190(.a(n3550), .b(n3556), .O(n3557));
  orx   g03191(.a(n3557), .b(n3555), .O(n3558));
  andx  g03192(.a(n3558), .b(n3553), .O(n3559));
  andx  g03193(.a(n3410), .b(n3312), .O(n3560));
  andx  g03194(.a(n3410), .b(n3407), .O(n3561));
  orx   g03195(.a(n3561), .b(n3560), .O(n3562));
  andx  g03196(.a(n3401), .b(n3153), .O(n3563));
  andx  g03197(.a(n3320), .b(n2668), .O(n3566));
  orx   g03198(.a(n3566), .b(n3322), .O(n3567));
  andx  g03199(.a(n3567), .b(n3319), .O(n3568));
  andx  g03200(.a(n2176), .b(n836), .O(n3569));
  invx  g03201(.a(n3569), .O(n3570));
  invx  g03202(.a(n3568), .O(n3572));
  andx  g03203(.a(n3569), .b(n3572), .O(n3573));
  orx   g03204(.a(n3573), .b(n830), .O(n3574));
  invx  g03205(.a(n3574), .O(n3575));
  andx  g03206(.a(n3575), .b(n2116), .O(n3576));
  andx  g03207(.a(n3574), .b(n2864), .O(n3577));
  orx   g03208(.a(n3577), .b(n3576), .O(n3578));
  andx  g03209(.a(n3337), .b(n3330), .O(n3579));
  orx   g03210(.a(n3579), .b(n3334), .O(n3580));
  invx  g03211(.a(n3580), .O(n3582));
  andx  g03212(.a(n605), .b(n3582), .O(n3585));
  invx  g03213(.a(n3585), .O(n3586));
  andx  g03214(.a(n3586), .b(n3578), .O(n3587));
  invx  g03215(.a(n3578), .O(n3588));
  andx  g03216(.a(n3585), .b(n3588), .O(n3589));
  orx   g03217(.a(n3589), .b(n3587), .O(n3590));
  invx  g03218(.a(n3590), .O(n3591));
  invx  g03219(.a(n3349), .O(n3593));
  andx  g03220(.a(n3349), .b(n3342), .O(n3596));
  orx   g03221(.a(n3596), .b(n560), .O(n3597));
  orx   g03222(.a(n3368), .b(n3591), .O(n3603));
  andx  g03223(.a(n3368), .b(n3591), .O(n3604));
  invx  g03224(.a(n3604), .O(n3605));
  andx  g03225(.a(n3605), .b(n3603), .O(n3606));
  andx  g03226(.a(n488), .b(n3359), .O(n3607));
  orx   g03227(.a(n3607), .b(n3361), .O(n3608));
  invx  g03228(.a(n3608), .O(n3612));
  andx  g03229(.a(n3612), .b(n3606), .O(n3614));
  invx  g03230(.a(n3603), .O(n3615));
  orx   g03231(.a(n3604), .b(n3615), .O(n3616));
  andx  g03232(.a(n3608), .b(n3616), .O(n3619));
  orx   g03233(.a(n3619), .b(n3614), .O(n3620));
  andx  g03234(.a(n3388), .b(n3620), .O(n3627));
  orx   g03235(.a(n3608), .b(n3616), .O(n3628));
  orx   g03236(.a(n3612), .b(n3606), .O(n3629));
  andx  g03237(.a(n3629), .b(n3628), .O(n3630));
  andx  g03238(.a(n3399), .b(n3630), .O(n3631));
  orx   g03239(.a(n3631), .b(n3627), .O(n3632));
  andx  g03240(.a(n3632), .b(n3563), .O(n3633));
  invx  g03241(.a(n3563), .O(n3634));
  orx   g03242(.a(n3399), .b(n3630), .O(n3635));
  orx   g03243(.a(n3388), .b(n3620), .O(n3636));
  andx  g03244(.a(n3636), .b(n3635), .O(n3637));
  andx  g03245(.a(n3637), .b(n3634), .O(n3638));
  orx   g03246(.a(n3638), .b(n3633), .O(n3639));
  andx  g03247(.a(n3639), .b(n3562), .O(n3640));
  orx   g03248(.a(n3637), .b(n3634), .O(n3641));
  orx   g03249(.a(n3632), .b(n3563), .O(n3642));
  andx  g03250(.a(n3642), .b(n3641), .O(n3643));
  andx  g03251(.a(n3643), .b(n3406), .O(n3644));
  orx   g03252(.a(n3644), .b(n3640), .O(n3645));
  andx  g03253(.a(n3645), .b(n299), .O(n3646));
  invx  g03254(.a(n3646), .O(n3647));
  andx  g03255(.a(n3647), .b(n3559), .O(n3648));
  invx  g03256(.a(n3559), .O(n3649));
  andx  g03257(.a(n3646), .b(n3649), .O(n3650));
  orx   g03258(.a(n3650), .b(n3648), .O(n3651));
  invx  g03259(.a(n3651), .O(n3652));
  andx  g03260(.a(n3652), .b(n3425), .O(n3653));
  andx  g03261(.a(n3651), .b(n3424), .O(n3654));
  orx   g03262(.a(n3654), .b(n3653), .O(n3655));
  invx  g03263(.a(n3655), .O(n3656));
  andx  g03264(.a(n3388), .b(n3630), .O(n3657));
  andx  g03265(.a(n3568), .b(n2864), .O(n3662));
  orx   g03266(.a(n3662), .b(n3570), .O(n3663));
  andx  g03267(.a(n3663), .b(n3567), .O(n3664));
  invx  g03268(.a(n3664), .O(n3668));
  orx   g03269(.a(n3668), .b(n830), .O(n3670));
  invx  g03270(.a(n3670), .O(n3671));
  orx   g03271(.a(n2333), .b(n3671), .O(n3674));
  andx  g03272(.a(n605), .b(n3588), .O(n3675));
  orx   g03273(.a(n3675), .b(n3580), .O(n3676));
  invx  g03274(.a(n3676), .O(n3678));
  andx  g03275(.a(n605), .b(n3678), .O(n3681));
  orx   g03276(.a(n3681), .b(n3674), .O(n3686));
  andx  g03277(.a(n2724), .b(n554), .O(n3687));
  invx  g03278(.a(n3687), .O(n3688));
  invx  g03279(.a(n3597), .O(n3689));
  andx  g03280(.a(n3689), .b(n3591), .O(n3690));
  andx  g03281(.a(n3597), .b(n3590), .O(n3691));
  invx  g03282(.a(n3691), .O(n3692));
  andx  g03283(.a(n3692), .b(n554), .O(n3693));
  orx   g03284(.a(n3693), .b(n3690), .O(n3694));
  andx  g03285(.a(n3694), .b(n3688), .O(n3695));
  invx  g03286(.a(n3694), .O(n3696));
  andx  g03287(.a(n3696), .b(n3687), .O(n3697));
  orx   g03288(.a(n3697), .b(n3695), .O(n3698));
  andx  g03289(.a(n3698), .b(n3686), .O(n3699));
  invx  g03290(.a(n3699), .O(n3700));
  orx   g03291(.a(n3698), .b(n3686), .O(n3701));
  andx  g03292(.a(n3701), .b(n3700), .O(n3702));
  orx   g03293(.a(n3702), .b(n3619), .O(n3703));
  invx  g03294(.a(n3703), .O(n3704));
  andx  g03295(.a(n3702), .b(n3619), .O(n3705));
  orx   g03296(.a(n3705), .b(n3704), .O(n3706));
  andx  g03297(.a(n3706), .b(n3657), .O(n3707));
  invx  g03298(.a(n3657), .O(n3708));
  invx  g03299(.a(n3705), .O(n3709));
  andx  g03300(.a(n3709), .b(n3703), .O(n3710));
  andx  g03301(.a(n3710), .b(n3708), .O(n3711));
  orx   g03302(.a(n3711), .b(n3707), .O(n3712));
  andx  g03303(.a(n3642), .b(n3562), .O(n3713));
  orx   g03304(.a(n3713), .b(n3633), .O(n3714));
  andx  g03305(.a(n3714), .b(n3712), .O(n3715));
  orx   g03306(.a(n3710), .b(n3708), .O(n3716));
  orx   g03307(.a(n3706), .b(n3657), .O(n3717));
  andx  g03308(.a(n3717), .b(n3716), .O(n3718));
  invx  g03309(.a(n3714), .O(n3719));
  andx  g03310(.a(n3719), .b(n3718), .O(n3720));
  orx   g03311(.a(n3720), .b(n3715), .O(n3721));
  invx  g03312(.a(n3511), .O(n3722));
  andx  g03313(.a(n3513), .b(n3473), .O(n3723));
  andx  g03314(.a(n3503), .b(n3512), .O(n3724));
  orx   g03315(.a(n3724), .b(n3723), .O(n3725));
  andx  g03316(.a(n3725), .b(n3722), .O(n3726));
  invx  g03317(.a(n3726), .O(n3727));
  orx   g03318(.a(n3725), .b(n3722), .O(n3728));
  andx  g03319(.a(n3728), .b(n3727), .O(n3729));
  invx  g03320(.a(n3729), .O(n3730));
  invx  g03321(.a(n3487), .O(n3731));
  andx  g03322(.a(n3501), .b(n3731), .O(n3732));
  invx  g03323(.a(n3732), .O(n3733));
  andx  g03324(.a(n3733), .b(n3499), .O(n3734));
  invx  g03325(.a(n3499), .O(n3735));
  andx  g03326(.a(n3732), .b(n3735), .O(n3736));
  orx   g03327(.a(n3736), .b(n3734), .O(n3737));
  andx  g03328(.a(n3210), .b(n338), .O(n3738));
  andx  g03329(.a(n3738), .b(n3737), .O(n3739));
  andx  g03330(.a(n3230), .b(n338), .O(n3740));
  andx  g03331(.a(n3258), .b(n338), .O(n3741));
  andx  g03332(.a(n1790), .b(n299), .O(n3742));
  andx  g03333(.a(n3742), .b(n3741), .O(n3743));
  andx  g03334(.a(n3743), .b(n3740), .O(n3744));
  invx  g03335(.a(n3475), .O(n3745));
  orx   g03336(.a(n3474), .b(n3241), .O(n3746));
  andx  g03337(.a(n3746), .b(n3745), .O(n3747));
  andx  g03338(.a(n3747), .b(n3740), .O(n3748));
  andx  g03339(.a(n3747), .b(n3743), .O(n3749));
  orx   g03340(.a(n3749), .b(n3748), .O(n3750));
  orx   g03341(.a(n3750), .b(n3744), .O(n3751));
  andx  g03342(.a(n3751), .b(n3221), .O(n3752));
  andx  g03343(.a(n3476), .b(n3745), .O(n3753));
  invx  g03344(.a(n3753), .O(n3754));
  orx   g03345(.a(n3476), .b(n3745), .O(n3755));
  andx  g03346(.a(n3755), .b(n3754), .O(n3756));
  andx  g03347(.a(n3756), .b(n3484), .O(n3757));
  invx  g03348(.a(n3757), .O(n3758));
  orx   g03349(.a(n3756), .b(n3484), .O(n3759));
  andx  g03350(.a(n3759), .b(n3758), .O(n3760));
  invx  g03351(.a(n3760), .O(n3761));
  andx  g03352(.a(n3221), .b(n338), .O(n3762));
  orx   g03353(.a(n3762), .b(n3751), .O(n3763));
  andx  g03354(.a(n3763), .b(n3761), .O(n3764));
  orx   g03355(.a(n3764), .b(n3752), .O(n3765));
  andx  g03356(.a(n3765), .b(n3737), .O(n3766));
  andx  g03357(.a(n3765), .b(n3738), .O(n3767));
  orx   g03358(.a(n3767), .b(n3766), .O(n3768));
  orx   g03359(.a(n3768), .b(n3739), .O(n3769));
  invx  g03360(.a(n3769), .O(n3770));
  andx  g03361(.a(n3770), .b(n3730), .O(n3771));
  andx  g03362(.a(n3284), .b(n338), .O(n3772));
  invx  g03363(.a(n3772), .O(n3773));
  orx   g03364(.a(n3773), .b(n3771), .O(n3774));
  andx  g03365(.a(n3769), .b(n3729), .O(n3775));
  invx  g03366(.a(n3775), .O(n3776));
  andx  g03367(.a(n3776), .b(n3774), .O(n3777));
  andx  g03368(.a(n3521), .b(n3517), .O(n3778));
  andx  g03369(.a(n3522), .b(n3516), .O(n3779));
  orx   g03370(.a(n3779), .b(n3778), .O(n3780));
  andx  g03371(.a(n3780), .b(n3471), .O(n3781));
  invx  g03372(.a(n3781), .O(n3782));
  orx   g03373(.a(n3780), .b(n3471), .O(n3783));
  andx  g03374(.a(n3783), .b(n3782), .O(n3784));
  andx  g03375(.a(n3966), .b(n3777), .O(n3786));
  andx  g03376(.a(n3180), .b(n338), .O(n3787));
  invx  g03377(.a(n3787), .O(n3788));
  andx  g03378(.a(n3788), .b(n3777), .O(n3789));
  andx  g03379(.a(n3788), .b(n3966), .O(n3790));
  orx   g03380(.a(n3790), .b(n3789), .O(n3791));
  orx   g03381(.a(n3791), .b(n3786), .O(n3792));
  invx  g03382(.a(n3792), .O(n3793));
  andx  g03383(.a(n3793), .b(n3429), .O(n3794));
  andx  g03384(.a(n3529), .b(n3525), .O(n3795));
  andx  g03385(.a(n3528), .b(n3524), .O(n3796));
  orx   g03386(.a(n3796), .b(n3795), .O(n3797));
  andx  g03387(.a(n3797), .b(n3530), .O(n3798));
  invx  g03388(.a(n3798), .O(n3799));
  orx   g03389(.a(n3797), .b(n3530), .O(n3800));
  andx  g03390(.a(n3800), .b(n3799), .O(n3801));
  invx  g03391(.a(n3801), .O(n3802));
  andx  g03392(.a(n3429), .b(n338), .O(n3803));
  orx   g03393(.a(n3803), .b(n3793), .O(n3804));
  andx  g03394(.a(n3804), .b(n3802), .O(n3805));
  orx   g03395(.a(n3805), .b(n3794), .O(n3806));
  andx  g03396(.a(n3806), .b(n3171), .O(n3807));
  andx  g03397(.a(n3537), .b(n3534), .O(n3808));
  andx  g03398(.a(n3538), .b(n3533), .O(n3809));
  orx   g03399(.a(n3809), .b(n3808), .O(n3810));
  invx  g03400(.a(n3810), .O(n3811));
  andx  g03401(.a(n3811), .b(n3539), .O(n3812));
  andx  g03402(.a(n3810), .b(n3454), .O(n3813));
  orx   g03403(.a(n3813), .b(n3812), .O(n3814));
  andx  g03404(.a(n3171), .b(n338), .O(n3815));
  orx   g03405(.a(n3815), .b(n3806), .O(n3816));
  andx  g03406(.a(n3816), .b(n3814), .O(n3817));
  orx   g03407(.a(n3817), .b(n3807), .O(n3818));
  andx  g03408(.a(n3818), .b(n3413), .O(n3819));
  andx  g03409(.a(n3547), .b(n3542), .O(n3820));
  andx  g03410(.a(n3546), .b(n3543), .O(n3821));
  orx   g03411(.a(n3821), .b(n3820), .O(n3822));
  invx  g03412(.a(n3822), .O(n3823));
  andx  g03413(.a(n3823), .b(n3445), .O(n3824));
  andx  g03414(.a(n3822), .b(n3446), .O(n3825));
  orx   g03415(.a(n3825), .b(n3824), .O(n3826));
  andx  g03416(.a(n3413), .b(n338), .O(n3827));
  orx   g03417(.a(n3827), .b(n3818), .O(n3828));
  andx  g03418(.a(n3828), .b(n3826), .O(n3829));
  orx   g03419(.a(n3829), .b(n3819), .O(n3830));
  andx  g03420(.a(n3830), .b(n3645), .O(n3831));
  andx  g03421(.a(n3555), .b(n3551), .O(n3832));
  andx  g03422(.a(n3554), .b(n3550), .O(n3833));
  orx   g03423(.a(n3833), .b(n3832), .O(n3834));
  andx  g03424(.a(n3834), .b(n3556), .O(n3835));
  invx  g03425(.a(n3835), .O(n3836));
  orx   g03426(.a(n3834), .b(n3556), .O(n3837));
  andx  g03427(.a(n3837), .b(n3836), .O(n3838));
  invx  g03428(.a(n3838), .O(n3839));
  andx  g03429(.a(n3645), .b(n338), .O(n3840));
  orx   g03430(.a(n3840), .b(n3830), .O(n3841));
  andx  g03431(.a(n3841), .b(n3839), .O(n3842));
  orx   g03432(.a(n3842), .b(n3831), .O(n3843));
  andx  g03433(.a(n3843), .b(n3721), .O(n3844));
  invx  g03434(.a(n3844), .O(n3845));
  andx  g03435(.a(n3721), .b(n338), .O(n3846));
  orx   g03436(.a(n3846), .b(n3843), .O(n3847));
  andx  g03437(.a(n3847), .b(n3845), .O(n3848));
  invx  g03438(.a(n3848), .O(n3849));
  andx  g03439(.a(n3849), .b(n3656), .O(n3850));
  andx  g03440(.a(n3848), .b(n3655), .O(n3851));
  orx   g03441(.a(n3851), .b(n3850), .O(n3852));
  invx  g03442(.a(n3831), .O(n3853));
  andx  g03443(.a(n3841), .b(n3853), .O(n3854));
  invx  g03444(.a(n3854), .O(n3855));
  andx  g03445(.a(n3855), .b(n3838), .O(n3856));
  andx  g03446(.a(n3854), .b(n3839), .O(n3857));
  orx   g03447(.a(n3857), .b(n3856), .O(n3858));
  invx  g03448(.a(n3826), .O(n3859));
  invx  g03449(.a(n3819), .O(n3860));
  andx  g03450(.a(n3828), .b(n3860), .O(n3861));
  invx  g03451(.a(n3861), .O(n3862));
  andx  g03452(.a(n3862), .b(n3859), .O(n3863));
  andx  g03453(.a(n3861), .b(n3826), .O(n3864));
  orx   g03454(.a(n3864), .b(n3863), .O(n3865));
  invx  g03455(.a(n3814), .O(n3866));
  invx  g03456(.a(n3807), .O(n3867));
  andx  g03457(.a(n3816), .b(n3867), .O(n3868));
  invx  g03458(.a(n3868), .O(n3869));
  andx  g03459(.a(n3869), .b(n3866), .O(n3870));
  andx  g03460(.a(n3868), .b(n3814), .O(n3871));
  orx   g03461(.a(n3871), .b(n3870), .O(n3872));
  invx  g03462(.a(n3794), .O(n3873));
  andx  g03463(.a(n3804), .b(n3873), .O(n3874));
  invx  g03464(.a(n3874), .O(n3875));
  andx  g03465(.a(n3875), .b(n3802), .O(n3876));
  andx  g03466(.a(n3874), .b(n3801), .O(n3877));
  orx   g03467(.a(n3877), .b(n3876), .O(n3878));
  invx  g03468(.a(n3878), .O(n3879));
  andx  g03469(.a(n3773), .b(n3769), .O(n3880));
  andx  g03470(.a(n3772), .b(n3770), .O(n3881));
  orx   g03471(.a(n3881), .b(n3880), .O(n3882));
  andx  g03472(.a(n3882), .b(n3730), .O(n3883));
  invx  g03473(.a(n3883), .O(n3884));
  orx   g03474(.a(n3882), .b(n3730), .O(n3885));
  andx  g03475(.a(n3885), .b(n3884), .O(n3886));
  invx  g03476(.a(n3886), .O(n3887));
  andx  g03477(.a(n3180), .b(n376), .O(n3888));
  andx  g03478(.a(n3888), .b(n3887), .O(n3889));
  invx  g03479(.a(n3889), .O(n3890));
  invx  g03480(.a(n3888), .O(n3891));
  andx  g03481(.a(n3891), .b(n3886), .O(n3892));
  andx  g03482(.a(n3210), .b(n376), .O(n3893));
  andx  g03483(.a(n3230), .b(n376), .O(n3894));
  invx  g03484(.a(n3742), .O(n3895));
  andx  g03485(.a(n3895), .b(n3741), .O(n3896));
  invx  g03486(.a(n3741), .O(n3897));
  andx  g03487(.a(n3742), .b(n3897), .O(n3898));
  orx   g03488(.a(n3898), .b(n3896), .O(n3899));
  andx  g03489(.a(n3899), .b(n3894), .O(n3900));
  andx  g03490(.a(n1790), .b(n338), .O(n3901));
  andx  g03491(.a(n3258), .b(n376), .O(n3902));
  andx  g03492(.a(n3902), .b(n3901), .O(n3903));
  andx  g03493(.a(n3903), .b(n3894), .O(n3904));
  andx  g03494(.a(n3903), .b(n3899), .O(n3905));
  orx   g03495(.a(n3905), .b(n3904), .O(n3906));
  orx   g03496(.a(n3906), .b(n3900), .O(n3907));
  andx  g03497(.a(n3907), .b(n3221), .O(n3908));
  invx  g03498(.a(n3743), .O(n3909));
  andx  g03499(.a(n3909), .b(n3740), .O(n3910));
  invx  g03500(.a(n3910), .O(n3911));
  orx   g03501(.a(n3909), .b(n3740), .O(n3912));
  andx  g03502(.a(n3912), .b(n3911), .O(n3913));
  andx  g03503(.a(n3913), .b(n3747), .O(n3914));
  invx  g03504(.a(n3914), .O(n3915));
  orx   g03505(.a(n3913), .b(n3747), .O(n3916));
  andx  g03506(.a(n3916), .b(n3915), .O(n3917));
  invx  g03507(.a(n3917), .O(n3918));
  andx  g03508(.a(n3221), .b(n376), .O(n3919));
  orx   g03509(.a(n3919), .b(n3907), .O(n3920));
  andx  g03510(.a(n3920), .b(n3918), .O(n3921));
  orx   g03511(.a(n3921), .b(n3908), .O(n3922));
  andx  g03512(.a(n3922), .b(n3893), .O(n3923));
  invx  g03513(.a(n3923), .O(n3924));
  invx  g03514(.a(n3752), .O(n3925));
  andx  g03515(.a(n3763), .b(n3925), .O(n3926));
  invx  g03516(.a(n3926), .O(n3927));
  andx  g03517(.a(n3927), .b(n3761), .O(n3928));
  andx  g03518(.a(n3926), .b(n3760), .O(n3929));
  orx   g03519(.a(n3929), .b(n3928), .O(n3930));
  invx  g03520(.a(n3930), .O(n3931));
  invx  g03521(.a(n3893), .O(n3932));
  invx  g03522(.a(n3922), .O(n3933));
  andx  g03523(.a(n3933), .b(n3932), .O(n3934));
  orx   g03524(.a(n3934), .b(n3931), .O(n3935));
  andx  g03525(.a(n3935), .b(n3924), .O(n3936));
  invx  g03526(.a(n3936), .O(n3937));
  andx  g03527(.a(n3937), .b(n3284), .O(n3938));
  invx  g03528(.a(n3738), .O(n3939));
  andx  g03529(.a(n3765), .b(n3939), .O(n3940));
  invx  g03530(.a(n3940), .O(n3941));
  orx   g03531(.a(n3765), .b(n3939), .O(n3942));
  andx  g03532(.a(n3942), .b(n3941), .O(n3943));
  invx  g03533(.a(n3943), .O(n3944));
  andx  g03534(.a(n3733), .b(n3735), .O(n3945));
  andx  g03535(.a(n3732), .b(n3499), .O(n3946));
  orx   g03536(.a(n3946), .b(n3945), .O(n3947));
  andx  g03537(.a(n3947), .b(n3944), .O(n3948));
  invx  g03538(.a(n3948), .O(n3949));
  orx   g03539(.a(n3947), .b(n3944), .O(n3950));
  andx  g03540(.a(n3950), .b(n3949), .O(n3951));
  invx  g03541(.a(n3951), .O(n3952));
  andx  g03542(.a(n3284), .b(n376), .O(n3953));
  orx   g03543(.a(n3953), .b(n3937), .O(n3954));
  andx  g03544(.a(n3954), .b(n3952), .O(n3955));
  orx   g03545(.a(n3955), .b(n3938), .O(n3956));
  invx  g03546(.a(n3956), .O(n3957));
  orx   g03547(.a(n3957), .b(n3892), .O(n3958));
  andx  g03548(.a(n3958), .b(n3890), .O(n3959));
  andx  g03549(.a(n3522), .b(n3517), .O(n3960));
  andx  g03550(.a(n3521), .b(n3516), .O(n3961));
  orx   g03551(.a(n3961), .b(n3960), .O(n3962));
  andx  g03552(.a(n3962), .b(n3471), .O(n3963));
  invx  g03553(.a(n3963), .O(n3964));
  orx   g03554(.a(n3962), .b(n3471), .O(n3965));
  andx  g03555(.a(n3965), .b(n3964), .O(n3966));
  invx  g03556(.a(n3777), .O(n3968));
  andx  g03557(.a(n3788), .b(n3968), .O(n3969));
  andx  g03558(.a(n3787), .b(n3777), .O(n3970));
  orx   g03559(.a(n3970), .b(n3969), .O(n3971));
  andx  g03560(.a(n3971), .b(n3784), .O(n3972));
  invx  g03561(.a(n3972), .O(n3973));
  orx   g03562(.a(n3971), .b(n3784), .O(n3974));
  andx  g03563(.a(n3974), .b(n3973), .O(n3975));
  invx  g03564(.a(n3975), .O(n3976));
  andx  g03565(.a(n3976), .b(n3959), .O(n3977));
  andx  g03566(.a(n3429), .b(n376), .O(n3978));
  invx  g03567(.a(n3978), .O(n3979));
  orx   g03568(.a(n3979), .b(n3977), .O(n3980));
  invx  g03569(.a(n3959), .O(n3981));
  andx  g03570(.a(n3975), .b(n3981), .O(n3982));
  invx  g03571(.a(n3982), .O(n3983));
  andx  g03572(.a(n3983), .b(n3980), .O(n3984));
  andx  g03573(.a(n3984), .b(n3879), .O(n3985));
  andx  g03574(.a(n3171), .b(n376), .O(n3986));
  invx  g03575(.a(n3986), .O(n3987));
  andx  g03576(.a(n3987), .b(n3879), .O(n3988));
  andx  g03577(.a(n3987), .b(n3984), .O(n3989));
  orx   g03578(.a(n3989), .b(n3988), .O(n3990));
  orx   g03579(.a(n3990), .b(n3985), .O(n3991));
  andx  g03580(.a(n3991), .b(n3872), .O(n3992));
  andx  g03581(.a(n3413), .b(n376), .O(n3993));
  invx  g03582(.a(n3993), .O(n3994));
  andx  g03583(.a(n3994), .b(n3872), .O(n3995));
  andx  g03584(.a(n3994), .b(n3991), .O(n3996));
  orx   g03585(.a(n3996), .b(n3995), .O(n3997));
  orx   g03586(.a(n3997), .b(n3992), .O(n3998));
  andx  g03587(.a(n3998), .b(n3865), .O(n3999));
  andx  g03588(.a(n3645), .b(n376), .O(n4000));
  invx  g03589(.a(n4000), .O(n4001));
  andx  g03590(.a(n4001), .b(n3865), .O(n4002));
  andx  g03591(.a(n4001), .b(n3998), .O(n4003));
  orx   g03592(.a(n4003), .b(n4002), .O(n4004));
  orx   g03593(.a(n4004), .b(n3999), .O(n4005));
  andx  g03594(.a(n4005), .b(n3858), .O(n4006));
  andx  g03595(.a(n3721), .b(n376), .O(n4007));
  invx  g03596(.a(n4007), .O(n4008));
  orx   g03597(.a(n4008), .b(n4006), .O(n4009));
  invx  g03598(.a(n3858), .O(n4010));
  invx  g03599(.a(n4005), .O(n4011));
  andx  g03600(.a(n4011), .b(n4010), .O(n4012));
  invx  g03601(.a(n4012), .O(n4013));
  andx  g03602(.a(n4013), .b(n4009), .O(n4014));
  invx  g03603(.a(n4014), .O(n4015));
  andx  g03604(.a(n2429), .b(n611), .O(n4039));
  invx  g03605(.a(n4039), .O(n4043));
  invx  g03606(.a(n3686), .O(n4044));
  andx  g03607(.a(n3694), .b(n4044), .O(n4047));
  invx  g03608(.a(n4047), .O(n4050));
  andx  g03609(.a(n4050), .b(n4043), .O(n4051));
  andx  g03610(.a(n4047), .b(n4039), .O(n4052));
  orx   g03611(.a(n4052), .b(n4051), .O(n4053));
  andx  g03612(.a(n3714), .b(n3717), .O(n4054));
  invx  g03613(.a(n3702), .O(n4055));
  andx  g03614(.a(n4055), .b(n3619), .O(n4056));
  orx   g03615(.a(n4056), .b(n3707), .O(n4057));
  orx   g03616(.a(n4057), .b(n4054), .O(n4058));
  andx  g03617(.a(n4058), .b(n4053), .O(n4059));
  invx  g03618(.a(n4059), .O(n4060));
  orx   g03619(.a(n4058), .b(n4053), .O(n4061));
  andx  g03620(.a(n4061), .b(n4060), .O(n4062));
  invx  g03621(.a(n4062), .O(n4063));
  andx  g03622(.a(n4063), .b(n376), .O(n4064));
  invx  g03623(.a(n4064), .O(n4065));
  andx  g03624(.a(n4065), .b(n4015), .O(n4066));
  andx  g03625(.a(n4064), .b(n4014), .O(n4067));
  orx   g03626(.a(n4067), .b(n4066), .O(n4068));
  andx  g03627(.a(n4068), .b(n3852), .O(n4069));
  invx  g03628(.a(n4069), .O(n4070));
  orx   g03629(.a(n4068), .b(n3852), .O(n4071));
  andx  g03630(.a(n4071), .b(n4070), .O(n4072));
  invx  g03631(.a(n4053), .O(n4073));
  andx  g03632(.a(n3642), .b(n3560), .O(n4074));
  orx   g03633(.a(n4074), .b(n3633), .O(n4075));
  andx  g03634(.a(n4075), .b(n3717), .O(n4076));
  orx   g03635(.a(n4076), .b(n4057), .O(n4077));
  andx  g03636(.a(n4077), .b(n4073), .O(n4078));
  andx  g03637(.a(n4073), .b(n3717), .O(n4079));
  andx  g03638(.a(n4079), .b(n3642), .O(n4080));
  andx  g03639(.a(n4080), .b(n3561), .O(n4081));
  orx   g03640(.a(n4081), .b(n4078), .O(n4082));
  invx  g03641(.a(n4082), .O(n4083));
  andx  g03642(.a(n830), .b(n2429), .O(n4100));
  andx  g03643(.a(n4100), .b(n611), .O(n4102));
  invx  g03644(.a(n4100), .O(n4103));
  andx  g03645(.a(n4103), .b(n605), .O(n4104));
  orx   g03646(.a(n4104), .b(n4102), .O(n4105));
  andx  g03647(.a(n4105), .b(n4052), .O(n4106));
  invx  g03648(.a(n4106), .O(n4107));
  orx   g03649(.a(n4105), .b(n4052), .O(n4108));
  andx  g03650(.a(n4108), .b(n4107), .O(n4109));
  invx  g03651(.a(n4109), .O(n4110));
  andx  g03652(.a(n4110), .b(n4083), .O(n4111));
  andx  g03653(.a(n4109), .b(n4082), .O(n4112));
  orx   g03654(.a(n4112), .b(n4111), .O(n4113));
  invx  g03655(.a(n4113), .O(n4114));
  andx  g03656(.a(n3956), .b(n3888), .O(n4115));
  andx  g03657(.a(n3957), .b(n3891), .O(n4116));
  orx   g03658(.a(n4116), .b(n4115), .O(n4117));
  invx  g03659(.a(n4117), .O(n4118));
  andx  g03660(.a(n4118), .b(n3887), .O(n4119));
  andx  g03661(.a(n4117), .b(n3886), .O(n4120));
  orx   g03662(.a(n4120), .b(n4119), .O(n4121));
  invx  g03663(.a(n4121), .O(n4122));
  invx  g03664(.a(n3938), .O(n4123));
  andx  g03665(.a(n3954), .b(n4123), .O(n4124));
  invx  g03666(.a(n4124), .O(n4125));
  andx  g03667(.a(n4125), .b(n3951), .O(n4126));
  andx  g03668(.a(n4124), .b(n3952), .O(n4127));
  orx   g03669(.a(n4127), .b(n4126), .O(n4128));
  invx  g03670(.a(n4128), .O(n4129));
  andx  g03671(.a(n3180), .b(n438), .O(n4130));
  andx  g03672(.a(n4130), .b(n4129), .O(n4131));
  invx  g03673(.a(n4131), .O(n4132));
  invx  g03674(.a(n4130), .O(n4133));
  andx  g03675(.a(n4133), .b(n4128), .O(n4134));
  andx  g03676(.a(n3933), .b(n3893), .O(n4135));
  andx  g03677(.a(n3922), .b(n3932), .O(n4136));
  orx   g03678(.a(n4136), .b(n4135), .O(n4137));
  andx  g03679(.a(n4137), .b(n3930), .O(n4138));
  invx  g03680(.a(n4138), .O(n4139));
  orx   g03681(.a(n4137), .b(n3930), .O(n4140));
  andx  g03682(.a(n4140), .b(n4139), .O(n4141));
  andx  g03683(.a(n3210), .b(n438), .O(n4142));
  andx  g03684(.a(n3230), .b(n438), .O(n4143));
  invx  g03685(.a(n3902), .O(n4144));
  andx  g03686(.a(n4144), .b(n3901), .O(n4145));
  invx  g03687(.a(n3901), .O(n4146));
  andx  g03688(.a(n3902), .b(n4146), .O(n4147));
  orx   g03689(.a(n4147), .b(n4145), .O(n4148));
  andx  g03690(.a(n4148), .b(n4143), .O(n4149));
  andx  g03691(.a(n1790), .b(n376), .O(n4150));
  andx  g03692(.a(n3258), .b(n438), .O(n4151));
  andx  g03693(.a(n4151), .b(n4150), .O(n4152));
  andx  g03694(.a(n4152), .b(n4143), .O(n4153));
  andx  g03695(.a(n4152), .b(n4148), .O(n4154));
  orx   g03696(.a(n4154), .b(n4153), .O(n4155));
  orx   g03697(.a(n4155), .b(n4149), .O(n4156));
  andx  g03698(.a(n4156), .b(n3221), .O(n4157));
  invx  g03699(.a(n3903), .O(n4158));
  andx  g03700(.a(n4158), .b(n3894), .O(n4159));
  invx  g03701(.a(n4159), .O(n4160));
  orx   g03702(.a(n4158), .b(n3894), .O(n4161));
  andx  g03703(.a(n4161), .b(n4160), .O(n4162));
  andx  g03704(.a(n3895), .b(n3897), .O(n4163));
  orx   g03705(.a(n4163), .b(n3743), .O(n4164));
  andx  g03706(.a(n4164), .b(n4162), .O(n4165));
  invx  g03707(.a(n4165), .O(n4166));
  orx   g03708(.a(n4164), .b(n4162), .O(n4167));
  andx  g03709(.a(n4167), .b(n4166), .O(n4168));
  andx  g03710(.a(n3221), .b(n438), .O(n4169));
  orx   g03711(.a(n4169), .b(n4156), .O(n4170));
  andx  g03712(.a(n4170), .b(n4168), .O(n4171));
  orx   g03713(.a(n4171), .b(n4157), .O(n4172));
  andx  g03714(.a(n4172), .b(n4142), .O(n4173));
  invx  g03715(.a(n4173), .O(n4174));
  invx  g03716(.a(n3908), .O(n4175));
  andx  g03717(.a(n3920), .b(n4175), .O(n4176));
  invx  g03718(.a(n4176), .O(n4177));
  andx  g03719(.a(n4177), .b(n3918), .O(n4178));
  andx  g03720(.a(n4176), .b(n3917), .O(n4179));
  orx   g03721(.a(n4179), .b(n4178), .O(n4180));
  invx  g03722(.a(n4180), .O(n4181));
  invx  g03723(.a(n4142), .O(n4182));
  invx  g03724(.a(n4172), .O(n4183));
  andx  g03725(.a(n4183), .b(n4182), .O(n4184));
  orx   g03726(.a(n4184), .b(n4181), .O(n4185));
  andx  g03727(.a(n4185), .b(n4174), .O(n4186));
  invx  g03728(.a(n4186), .O(n4187));
  andx  g03729(.a(n4187), .b(n4141), .O(n4188));
  invx  g03730(.a(n4188), .O(n4189));
  invx  g03731(.a(n4141), .O(n4190));
  andx  g03732(.a(n4186), .b(n4190), .O(n4191));
  andx  g03733(.a(n3284), .b(n438), .O(n4192));
  invx  g03734(.a(n4192), .O(n4193));
  orx   g03735(.a(n4193), .b(n4191), .O(n4194));
  andx  g03736(.a(n4194), .b(n4189), .O(n4195));
  orx   g03737(.a(n4195), .b(n4134), .O(n4196));
  andx  g03738(.a(n4196), .b(n4132), .O(n4197));
  invx  g03739(.a(n4197), .O(n4198));
  andx  g03740(.a(n4198), .b(n4122), .O(n4199));
  invx  g03741(.a(n4199), .O(n4200));
  andx  g03742(.a(n4197), .b(n4121), .O(n4201));
  andx  g03743(.a(n3429), .b(n438), .O(n4202));
  invx  g03744(.a(n4202), .O(n4203));
  orx   g03745(.a(n4203), .b(n4201), .O(n4204));
  andx  g03746(.a(n4204), .b(n4200), .O(n4205));
  invx  g03747(.a(n4205), .O(n4206));
  andx  g03748(.a(n4206), .b(n3171), .O(n4207));
  andx  g03749(.a(n3979), .b(n3981), .O(n4208));
  andx  g03750(.a(n3978), .b(n3959), .O(n4209));
  orx   g03751(.a(n4209), .b(n4208), .O(n4210));
  andx  g03752(.a(n4210), .b(n3976), .O(n4211));
  invx  g03753(.a(n4211), .O(n4212));
  orx   g03754(.a(n4210), .b(n3976), .O(n4213));
  andx  g03755(.a(n4213), .b(n4212), .O(n4214));
  invx  g03756(.a(n4214), .O(n4215));
  andx  g03757(.a(n3171), .b(n438), .O(n4216));
  orx   g03758(.a(n4216), .b(n4206), .O(n4217));
  andx  g03759(.a(n4217), .b(n4215), .O(n4218));
  orx   g03760(.a(n4218), .b(n4207), .O(n4219));
  andx  g03761(.a(n4219), .b(n3413), .O(n4220));
  invx  g03762(.a(n3984), .O(n4221));
  andx  g03763(.a(n3987), .b(n4221), .O(n4222));
  andx  g03764(.a(n3986), .b(n3984), .O(n4223));
  orx   g03765(.a(n4223), .b(n4222), .O(n4224));
  andx  g03766(.a(n4224), .b(n3878), .O(n4225));
  invx  g03767(.a(n4225), .O(n4226));
  orx   g03768(.a(n4224), .b(n3878), .O(n4227));
  andx  g03769(.a(n4227), .b(n4226), .O(n4228));
  andx  g03770(.a(n3413), .b(n438), .O(n4229));
  orx   g03771(.a(n4229), .b(n4219), .O(n4230));
  andx  g03772(.a(n4230), .b(n4228), .O(n4231));
  orx   g03773(.a(n4231), .b(n4220), .O(n4232));
  andx  g03774(.a(n4232), .b(n3645), .O(n4233));
  invx  g03775(.a(n3872), .O(n4234));
  invx  g03776(.a(n3996), .O(n4235));
  orx   g03777(.a(n3994), .b(n3991), .O(n4236));
  andx  g03778(.a(n4236), .b(n4235), .O(n4237));
  andx  g03779(.a(n4237), .b(n4234), .O(n4238));
  invx  g03780(.a(n4238), .O(n4239));
  orx   g03781(.a(n4237), .b(n4234), .O(n4240));
  andx  g03782(.a(n4240), .b(n4239), .O(n4241));
  andx  g03783(.a(n3645), .b(n438), .O(n4242));
  orx   g03784(.a(n4242), .b(n4232), .O(n4243));
  andx  g03785(.a(n4243), .b(n4241), .O(n4244));
  orx   g03786(.a(n4244), .b(n4233), .O(n4245));
  andx  g03787(.a(n4245), .b(n3721), .O(n4246));
  invx  g03788(.a(n3865), .O(n4247));
  invx  g03789(.a(n4003), .O(n4248));
  orx   g03790(.a(n4001), .b(n3998), .O(n4249));
  andx  g03791(.a(n4249), .b(n4248), .O(n4250));
  andx  g03792(.a(n4250), .b(n4247), .O(n4251));
  invx  g03793(.a(n4251), .O(n4252));
  orx   g03794(.a(n4250), .b(n4247), .O(n4253));
  andx  g03795(.a(n4253), .b(n4252), .O(n4254));
  andx  g03796(.a(n3721), .b(n438), .O(n4255));
  orx   g03797(.a(n4255), .b(n4245), .O(n4256));
  andx  g03798(.a(n4256), .b(n4254), .O(n4257));
  orx   g03799(.a(n4257), .b(n4246), .O(n4258));
  andx  g03800(.a(n4258), .b(n4063), .O(n4259));
  andx  g03801(.a(n4007), .b(n4011), .O(n4260));
  andx  g03802(.a(n4008), .b(n4005), .O(n4261));
  orx   g03803(.a(n4261), .b(n4260), .O(n4262));
  invx  g03804(.a(n4262), .O(n4263));
  andx  g03805(.a(n4263), .b(n4010), .O(n4264));
  andx  g03806(.a(n4262), .b(n3858), .O(n4265));
  orx   g03807(.a(n4265), .b(n4264), .O(n4266));
  invx  g03808(.a(n4266), .O(n4267));
  andx  g03809(.a(n4063), .b(n438), .O(n4268));
  orx   g03810(.a(n4268), .b(n4258), .O(n4269));
  andx  g03811(.a(n4269), .b(n4267), .O(n4270));
  orx   g03812(.a(n4270), .b(n4259), .O(n4271));
  andx  g03813(.a(n4271), .b(n4114), .O(n4272));
  invx  g03814(.a(n4272), .O(n4273));
  andx  g03815(.a(n4114), .b(n438), .O(n4274));
  orx   g03816(.a(n4274), .b(n4271), .O(n4275));
  andx  g03817(.a(n4275), .b(n4273), .O(n4276));
  invx  g03818(.a(n4276), .O(n4277));
  andx  g03819(.a(n4277), .b(n4072), .O(n4278));
  invx  g03820(.a(n4072), .O(n4279));
  andx  g03821(.a(n4276), .b(n4279), .O(n4280));
  orx   g03822(.a(n4280), .b(n4278), .O(n4281));
  invx  g03823(.a(n4259), .O(n4282));
  andx  g03824(.a(n4269), .b(n4282), .O(n4283));
  invx  g03825(.a(n4283), .O(n4284));
  andx  g03826(.a(n4284), .b(n4266), .O(n4285));
  andx  g03827(.a(n4283), .b(n4267), .O(n4286));
  orx   g03828(.a(n4286), .b(n4285), .O(n4287));
  invx  g03829(.a(n4287), .O(n4288));
  invx  g03830(.a(n4241), .O(n4289));
  invx  g03831(.a(n4233), .O(n4290));
  andx  g03832(.a(n4243), .b(n4290), .O(n4291));
  invx  g03833(.a(n4291), .O(n4292));
  andx  g03834(.a(n4292), .b(n4289), .O(n4293));
  andx  g03835(.a(n4291), .b(n4241), .O(n4294));
  orx   g03836(.a(n4294), .b(n4293), .O(n4295));
  invx  g03837(.a(n4295), .O(n4296));
  invx  g03838(.a(n4228), .O(n4297));
  invx  g03839(.a(n4220), .O(n4298));
  andx  g03840(.a(n4230), .b(n4298), .O(n4299));
  invx  g03841(.a(n4299), .O(n4300));
  andx  g03842(.a(n4300), .b(n4297), .O(n4301));
  andx  g03843(.a(n4299), .b(n4228), .O(n4302));
  orx   g03844(.a(n4302), .b(n4301), .O(n4303));
  invx  g03845(.a(n4303), .O(n4304));
  invx  g03846(.a(n4207), .O(n4305));
  andx  g03847(.a(n4217), .b(n4305), .O(n4306));
  orx   g03848(.a(n4306), .b(n4215), .O(n4307));
  andx  g03849(.a(n4306), .b(n4215), .O(n4308));
  invx  g03850(.a(n4308), .O(n4309));
  andx  g03851(.a(n4309), .b(n4307), .O(n4310));
  invx  g03852(.a(n4310), .O(n4311));
  andx  g03853(.a(n4195), .b(n4133), .O(n4312));
  invx  g03854(.a(n4312), .O(n4313));
  orx   g03855(.a(n4195), .b(n4133), .O(n4314));
  andx  g03856(.a(n4314), .b(n4313), .O(n4315));
  andx  g03857(.a(n4315), .b(n4129), .O(n4316));
  invx  g03858(.a(n4316), .O(n4317));
  orx   g03859(.a(n4315), .b(n4129), .O(n4318));
  andx  g03860(.a(n4318), .b(n4317), .O(n4319));
  invx  g03861(.a(n4157), .O(n4320));
  andx  g03862(.a(n4170), .b(n4320), .O(n4321));
  invx  g03863(.a(n4321), .O(n4322));
  andx  g03864(.a(n4322), .b(n4168), .O(n4323));
  invx  g03865(.a(n4323), .O(n4324));
  orx   g03866(.a(n4322), .b(n4168), .O(n4325));
  andx  g03867(.a(n4325), .b(n4324), .O(n4326));
  invx  g03868(.a(n4326), .O(n4327));
  andx  g03869(.a(n3230), .b(n252), .O(n4328));
  invx  g03870(.a(n4151), .O(n4329));
  andx  g03871(.a(n4329), .b(n4150), .O(n4330));
  invx  g03872(.a(n4150), .O(n4331));
  andx  g03873(.a(n4151), .b(n4331), .O(n4332));
  orx   g03874(.a(n4332), .b(n4330), .O(n4333));
  andx  g03875(.a(n4333), .b(n4328), .O(n4334));
  andx  g03876(.a(n1790), .b(n438), .O(n4335));
  andx  g03877(.a(n3258), .b(n252), .O(n4336));
  andx  g03878(.a(n4336), .b(n4335), .O(n4337));
  andx  g03879(.a(n4337), .b(n4328), .O(n4338));
  andx  g03880(.a(n4337), .b(n4333), .O(n4339));
  orx   g03881(.a(n4339), .b(n4338), .O(n4340));
  orx   g03882(.a(n4340), .b(n4334), .O(n4341));
  andx  g03883(.a(n4341), .b(n3221), .O(n4342));
  andx  g03884(.a(n4144), .b(n4146), .O(n4343));
  orx   g03885(.a(n4343), .b(n3903), .O(n4344));
  invx  g03886(.a(n4153), .O(n4345));
  orx   g03887(.a(n4152), .b(n4143), .O(n4346));
  andx  g03888(.a(n4346), .b(n4345), .O(n4347));
  invx  g03889(.a(n4347), .O(n4348));
  andx  g03890(.a(n4348), .b(n4344), .O(n4349));
  invx  g03891(.a(n4349), .O(n4350));
  orx   g03892(.a(n4348), .b(n4344), .O(n4351));
  andx  g03893(.a(n4351), .b(n4350), .O(n4352));
  andx  g03894(.a(n3221), .b(n252), .O(n4353));
  orx   g03895(.a(n4353), .b(n4341), .O(n4354));
  andx  g03896(.a(n4354), .b(n4352), .O(n4355));
  orx   g03897(.a(n4355), .b(n4342), .O(n4356));
  andx  g03898(.a(n4356), .b(n4327), .O(n4357));
  invx  g03899(.a(n4357), .O(n4358));
  andx  g03900(.a(n3210), .b(n252), .O(n4359));
  invx  g03901(.a(n4359), .O(n4360));
  invx  g03902(.a(n4356), .O(n4361));
  andx  g03903(.a(n4361), .b(n4326), .O(n4362));
  orx   g03904(.a(n4362), .b(n4360), .O(n4363));
  andx  g03905(.a(n4363), .b(n4358), .O(n4364));
  andx  g03906(.a(n4172), .b(n4182), .O(n4365));
  andx  g03907(.a(n4183), .b(n4142), .O(n4366));
  orx   g03908(.a(n4366), .b(n4365), .O(n4367));
  andx  g03909(.a(n4367), .b(n4181), .O(n4368));
  invx  g03910(.a(n4368), .O(n4369));
  orx   g03911(.a(n4367), .b(n4181), .O(n4370));
  andx  g03912(.a(n4370), .b(n4369), .O(n4371));
  andx  g03913(.a(n4371), .b(n4364), .O(n4372));
  andx  g03914(.a(n3284), .b(n252), .O(n4373));
  invx  g03915(.a(n4373), .O(n4374));
  orx   g03916(.a(n4374), .b(n4372), .O(n4375));
  invx  g03917(.a(n4364), .O(n4376));
  invx  g03918(.a(n4371), .O(n4377));
  andx  g03919(.a(n4377), .b(n4376), .O(n4378));
  invx  g03920(.a(n4378), .O(n4379));
  andx  g03921(.a(n4379), .b(n4375), .O(n4380));
  andx  g03922(.a(n4192), .b(n4186), .O(n4381));
  andx  g03923(.a(n4193), .b(n4187), .O(n4382));
  orx   g03924(.a(n4382), .b(n4381), .O(n4383));
  andx  g03925(.a(n4536), .b(n4190), .O(n4385));
  andx  g03926(.a(n4383), .b(n4141), .O(n4386));
  orx   g03927(.a(n4386), .b(n4385), .O(n4387));
  andx  g03928(.a(n4387), .b(n4380), .O(n4388));
  andx  g03929(.a(n3180), .b(n252), .O(n4389));
  invx  g03930(.a(n4389), .O(n4390));
  andx  g03931(.a(n4390), .b(n4380), .O(n4391));
  andx  g03932(.a(n4390), .b(n4387), .O(n4392));
  orx   g03933(.a(n4392), .b(n4391), .O(n4393));
  orx   g03934(.a(n4393), .b(n4388), .O(n4394));
  invx  g03935(.a(n4394), .O(n4395));
  andx  g03936(.a(n4395), .b(n4319), .O(n4396));
  andx  g03937(.a(n3429), .b(n252), .O(n4397));
  orx   g03938(.a(n4395), .b(n4319), .O(n4398));
  andx  g03939(.a(n4398), .b(n4397), .O(n4399));
  orx   g03940(.a(n4399), .b(n4396), .O(n4400));
  invx  g03941(.a(n4400), .O(n4401));
  andx  g03942(.a(n3171), .b(n252), .O(n4402));
  invx  g03943(.a(n4402), .O(n4403));
  andx  g03944(.a(n4203), .b(n4198), .O(n4404));
  andx  g03945(.a(n4202), .b(n4197), .O(n4405));
  orx   g03946(.a(n4405), .b(n4404), .O(n4406));
  andx  g03947(.a(n4406), .b(n4121), .O(n4407));
  invx  g03948(.a(n4407), .O(n4408));
  orx   g03949(.a(n4406), .b(n4121), .O(n4409));
  andx  g03950(.a(n4409), .b(n4408), .O(n4410));
  andx  g03951(.a(n4410), .b(n4403), .O(n4411));
  orx   g03952(.a(n4411), .b(n4401), .O(n4412));
  invx  g03953(.a(n4410), .O(n4413));
  andx  g03954(.a(n4413), .b(n4402), .O(n4414));
  invx  g03955(.a(n4414), .O(n4415));
  andx  g03956(.a(n4415), .b(n4412), .O(n4416));
  andx  g03957(.a(n4416), .b(n4311), .O(n4417));
  andx  g03958(.a(n3413), .b(n252), .O(n4418));
  invx  g03959(.a(n4418), .O(n4419));
  andx  g03960(.a(n4419), .b(n4311), .O(n4420));
  andx  g03961(.a(n4419), .b(n4416), .O(n4421));
  orx   g03962(.a(n4421), .b(n4420), .O(n4422));
  orx   g03963(.a(n4422), .b(n4417), .O(n4423));
  invx  g03964(.a(n4423), .O(n4424));
  andx  g03965(.a(n4424), .b(n4304), .O(n4425));
  invx  g03966(.a(n4425), .O(n4426));
  andx  g03967(.a(n3645), .b(n252), .O(n4427));
  invx  g03968(.a(n4427), .O(n4428));
  andx  g03969(.a(n4423), .b(n4303), .O(n4429));
  orx   g03970(.a(n4429), .b(n4428), .O(n4430));
  andx  g03971(.a(n4430), .b(n4426), .O(n4431));
  invx  g03972(.a(n4431), .O(n4432));
  andx  g03973(.a(n4432), .b(n4296), .O(n4433));
  invx  g03974(.a(n4433), .O(n4434));
  andx  g03975(.a(n3721), .b(n252), .O(n4435));
  invx  g03976(.a(n4435), .O(n4436));
  andx  g03977(.a(n4431), .b(n4295), .O(n4437));
  orx   g03978(.a(n4437), .b(n4436), .O(n4438));
  andx  g03979(.a(n4438), .b(n4434), .O(n4439));
  invx  g03980(.a(n4254), .O(n4440));
  invx  g03981(.a(n4246), .O(n4441));
  andx  g03982(.a(n4256), .b(n4441), .O(n4442));
  invx  g03983(.a(n4442), .O(n4443));
  andx  g03984(.a(n4443), .b(n4440), .O(n4444));
  andx  g03985(.a(n4442), .b(n4254), .O(n4445));
  orx   g03986(.a(n4445), .b(n4444), .O(n4446));
  andx  g03987(.a(n4446), .b(n4439), .O(n4447));
  andx  g03988(.a(n4063), .b(n252), .O(n4448));
  invx  g03989(.a(n4448), .O(n4449));
  orx   g03990(.a(n4449), .b(n4447), .O(n4450));
  invx  g03991(.a(n4439), .O(n4451));
  invx  g03992(.a(n4446), .O(n4452));
  andx  g03993(.a(n4452), .b(n4451), .O(n4453));
  invx  g03994(.a(n4453), .O(n4454));
  andx  g03995(.a(n4454), .b(n4450), .O(n4455));
  invx  g03996(.a(n4455), .O(n4456));
  andx  g03997(.a(n4456), .b(n4288), .O(n4457));
  invx  g03998(.a(n4457), .O(n4458));
  andx  g03999(.a(n4455), .b(n4287), .O(n4459));
  andx  g04000(.a(n4114), .b(n252), .O(n4460));
  invx  g04001(.a(n4460), .O(n4461));
  orx   g04002(.a(n4461), .b(n4459), .O(n4462));
  andx  g04003(.a(n4462), .b(n4458), .O(n4463));
  invx  g04004(.a(n4463), .O(n4464));
  invx  g04005(.a(n2074), .O(n4466));
  orx   g04006(.a(n4112), .b(n4106), .O(n4468));
  invx  g04007(.a(n4468), .O(n4469));
  andx  g04008(.a(n4469), .b(n4466), .O(n4470));
  orx   g04009(.a(n1136), .b(n836), .O(n4485));
  invx  g04010(.a(n4485), .O(n4486));
  andx  g04011(.a(n4486), .b(n4470), .O(n4487));
  invx  g04012(.a(n4487), .O(n4488));
  orx   g04013(.a(n4486), .b(n4470), .O(n4489));
  andx  g04014(.a(n4489), .b(n4488), .O(n4490));
  andx  g04015(.a(n4490), .b(n252), .O(n4491));
  invx  g04016(.a(n4491), .O(n4492));
  andx  g04017(.a(n4492), .b(n4464), .O(n4493));
  andx  g04018(.a(n4491), .b(n4463), .O(n4494));
  orx   g04019(.a(n4494), .b(n4493), .O(n4495));
  andx  g04020(.a(n4495), .b(n4281), .O(n4496));
  invx  g04021(.a(n4496), .O(n4497));
  orx   g04022(.a(n4495), .b(n4281), .O(n4498));
  andx  g04023(.a(n4498), .b(n4497), .O(n4499));
  orx   g04024(.a(n3643), .b(n3406), .O(n4507));
  orx   g04025(.a(n3639), .b(n3562), .O(n4508));
  andx  g04026(.a(n4508), .b(n4507), .O(n4509));
  andx  g04027(.a(n4403), .b(n4400), .O(n4510));
  invx  g04028(.a(n4510), .O(n4511));
  orx   g04029(.a(n4403), .b(n4400), .O(n4512));
  andx  g04030(.a(n4512), .b(n4511), .O(n4513));
  invx  g04031(.a(n4513), .O(n4514));
  andx  g04032(.a(n4514), .b(n4413), .O(n4515));
  andx  g04033(.a(n4513), .b(n4410), .O(n4516));
  orx   g04034(.a(n4516), .b(n4515), .O(n4517));
  invx  g04035(.a(n4517), .O(n4518));
  invx  g04036(.a(n4319), .O(n4519));
  andx  g04037(.a(n4397), .b(n4395), .O(n4520));
  invx  g04038(.a(n4520), .O(n4521));
  orx   g04039(.a(n4397), .b(n4395), .O(n4522));
  andx  g04040(.a(n4522), .b(n4521), .O(n4523));
  andx  g04041(.a(n4523), .b(n4519), .O(n4524));
  invx  g04042(.a(n4524), .O(n4525));
  orx   g04043(.a(n4523), .b(n4519), .O(n4526));
  andx  g04044(.a(n4526), .b(n4525), .O(n4527));
  invx  g04045(.a(n4527), .O(n4528));
  andx  g04046(.a(n3171), .b(n214), .O(n4529));
  andx  g04047(.a(n4529), .b(n4528), .O(n4530));
  invx  g04048(.a(n4530), .O(n4531));
  invx  g04049(.a(n4529), .O(n4532));
  andx  g04050(.a(n4532), .b(n4527), .O(n4533));
  andx  g04051(.a(n4193), .b(n4186), .O(n4534));
  andx  g04052(.a(n4192), .b(n4187), .O(n4535));
  orx   g04053(.a(n4535), .b(n4534), .O(n4536));
  andx  g04054(.a(n4383), .b(n4190), .O(n4538));
  andx  g04055(.a(n4536), .b(n4141), .O(n4539));
  orx   g04056(.a(n4539), .b(n4538), .O(n4540));
  invx  g04057(.a(n4391), .O(n4541));
  orx   g04058(.a(n4390), .b(n4380), .O(n4542));
  andx  g04059(.a(n4542), .b(n4541), .O(n4543));
  andx  g04060(.a(n4543), .b(n4540), .O(n4544));
  invx  g04061(.a(n4544), .O(n4545));
  orx   g04062(.a(n4543), .b(n4540), .O(n4546));
  andx  g04063(.a(n4546), .b(n4545), .O(n4547));
  orx   g04064(.a(n4373), .b(n4364), .O(n4548));
  andx  g04065(.a(n4373), .b(n4364), .O(n4549));
  invx  g04066(.a(n4549), .O(n4550));
  andx  g04067(.a(n4550), .b(n4548), .O(n4551));
  invx  g04068(.a(n4551), .O(n4552));
  andx  g04069(.a(n4552), .b(n4377), .O(n4553));
  andx  g04070(.a(n4551), .b(n4371), .O(n4554));
  orx   g04071(.a(n4554), .b(n4553), .O(n4555));
  invx  g04072(.a(n4555), .O(n4556));
  orx   g04073(.a(n4359), .b(n4356), .O(n4557));
  andx  g04074(.a(n4359), .b(n4356), .O(n4558));
  invx  g04075(.a(n4558), .O(n4559));
  andx  g04076(.a(n4559), .b(n4557), .O(n4560));
  andx  g04077(.a(n4560), .b(n4326), .O(n4561));
  invx  g04078(.a(n4561), .O(n4562));
  orx   g04079(.a(n4560), .b(n4326), .O(n4563));
  andx  g04080(.a(n4563), .b(n4562), .O(n4564));
  invx  g04081(.a(n4564), .O(n4565));
  invx  g04082(.a(n4342), .O(n4566));
  andx  g04083(.a(n4354), .b(n4566), .O(n4567));
  invx  g04084(.a(n4567), .O(n4568));
  andx  g04085(.a(n4568), .b(n4352), .O(n4569));
  invx  g04086(.a(n4569), .O(n4570));
  orx   g04087(.a(n4568), .b(n4352), .O(n4571));
  andx  g04088(.a(n4571), .b(n4570), .O(n4572));
  invx  g04089(.a(n4572), .O(n4573));
  andx  g04090(.a(n3230), .b(n214), .O(n4574));
  invx  g04091(.a(n4336), .O(n4575));
  andx  g04092(.a(n4575), .b(n4335), .O(n4576));
  invx  g04093(.a(n4335), .O(n4577));
  andx  g04094(.a(n4336), .b(n4577), .O(n4578));
  orx   g04095(.a(n4578), .b(n4576), .O(n4579));
  andx  g04096(.a(n4579), .b(n4574), .O(n4580));
  andx  g04097(.a(n1790), .b(n252), .O(n4581));
  andx  g04098(.a(n3258), .b(n214), .O(n4582));
  andx  g04099(.a(n4582), .b(n4581), .O(n4583));
  andx  g04100(.a(n4583), .b(n4574), .O(n4584));
  andx  g04101(.a(n4583), .b(n4579), .O(n4585));
  orx   g04102(.a(n4585), .b(n4584), .O(n4586));
  orx   g04103(.a(n4586), .b(n4580), .O(n4587));
  andx  g04104(.a(n4587), .b(n3221), .O(n4588));
  invx  g04105(.a(n4337), .O(n4589));
  andx  g04106(.a(n4589), .b(n4328), .O(n4590));
  invx  g04107(.a(n4590), .O(n4591));
  orx   g04108(.a(n4589), .b(n4328), .O(n4592));
  andx  g04109(.a(n4592), .b(n4591), .O(n4593));
  andx  g04110(.a(n4329), .b(n4331), .O(n4594));
  orx   g04111(.a(n4594), .b(n4152), .O(n4595));
  andx  g04112(.a(n4595), .b(n4593), .O(n4596));
  invx  g04113(.a(n4596), .O(n4597));
  orx   g04114(.a(n4595), .b(n4593), .O(n4598));
  andx  g04115(.a(n4598), .b(n4597), .O(n4599));
  andx  g04116(.a(n3221), .b(n214), .O(n4600));
  orx   g04117(.a(n4600), .b(n4587), .O(n4601));
  andx  g04118(.a(n4601), .b(n4599), .O(n4602));
  orx   g04119(.a(n4602), .b(n4588), .O(n4603));
  andx  g04120(.a(n4603), .b(n4573), .O(n4604));
  invx  g04121(.a(n4604), .O(n4605));
  andx  g04122(.a(n3210), .b(n214), .O(n4606));
  invx  g04123(.a(n4606), .O(n4607));
  invx  g04124(.a(n4603), .O(n4608));
  andx  g04125(.a(n4608), .b(n4572), .O(n4609));
  orx   g04126(.a(n4609), .b(n4607), .O(n4610));
  andx  g04127(.a(n4610), .b(n4605), .O(n4611));
  invx  g04128(.a(n4611), .O(n4612));
  andx  g04129(.a(n4612), .b(n4565), .O(n4613));
  invx  g04130(.a(n4613), .O(n4614));
  andx  g04131(.a(n4611), .b(n4564), .O(n4615));
  andx  g04132(.a(n3284), .b(n214), .O(n4616));
  invx  g04133(.a(n4616), .O(n4617));
  orx   g04134(.a(n4617), .b(n4615), .O(n4618));
  andx  g04135(.a(n4618), .b(n4614), .O(n4619));
  invx  g04136(.a(n4619), .O(n4620));
  andx  g04137(.a(n4620), .b(n4556), .O(n4621));
  invx  g04138(.a(n4621), .O(n4622));
  andx  g04139(.a(n3180), .b(n214), .O(n4623));
  invx  g04140(.a(n4623), .O(n4624));
  andx  g04141(.a(n4619), .b(n4555), .O(n4625));
  orx   g04142(.a(n4625), .b(n4624), .O(n4626));
  andx  g04143(.a(n4626), .b(n4622), .O(n4627));
  invx  g04144(.a(n4627), .O(n4628));
  andx  g04145(.a(n4628), .b(n4547), .O(n4629));
  invx  g04146(.a(n4629), .O(n4630));
  andx  g04147(.a(n3429), .b(n214), .O(n4631));
  invx  g04148(.a(n4631), .O(n4632));
  invx  g04149(.a(n4547), .O(n4633));
  andx  g04150(.a(n4627), .b(n4633), .O(n4634));
  orx   g04151(.a(n4634), .b(n4632), .O(n4635));
  andx  g04152(.a(n4635), .b(n4630), .O(n4636));
  orx   g04153(.a(n4636), .b(n4533), .O(n4637));
  andx  g04154(.a(n4637), .b(n4531), .O(n4638));
  invx  g04155(.a(n4638), .O(n4639));
  andx  g04156(.a(n4639), .b(n4518), .O(n4640));
  invx  g04157(.a(n4640), .O(n4641));
  andx  g04158(.a(n3413), .b(n214), .O(n4642));
  invx  g04159(.a(n4642), .O(n4643));
  andx  g04160(.a(n4638), .b(n4517), .O(n4644));
  orx   g04161(.a(n4644), .b(n4643), .O(n4645));
  andx  g04162(.a(n4645), .b(n4641), .O(n4646));
  orx   g04163(.a(n4646), .b(n4509), .O(n4647));
  invx  g04164(.a(n4647), .O(n4648));
  invx  g04165(.a(n4421), .O(n4649));
  orx   g04166(.a(n4419), .b(n4416), .O(n4650));
  andx  g04167(.a(n4650), .b(n4649), .O(n4651));
  andx  g04168(.a(n4651), .b(n4310), .O(n4652));
  invx  g04169(.a(n4652), .O(n4653));
  orx   g04170(.a(n4651), .b(n4310), .O(n4654));
  andx  g04171(.a(n4654), .b(n4653), .O(n4655));
  andx  g04172(.a(n3645), .b(n214), .O(n4656));
  invx  g04173(.a(n4656), .O(n4657));
  andx  g04174(.a(n4657), .b(n4646), .O(n4658));
  invx  g04175(.a(n4658), .O(n4659));
  andx  g04176(.a(n4659), .b(n4655), .O(n4660));
  orx   g04177(.a(n4660), .b(n4648), .O(n4661));
  andx  g04178(.a(n4661), .b(n3721), .O(n4662));
  andx  g04179(.a(n4427), .b(n4424), .O(n4663));
  andx  g04180(.a(n4428), .b(n4423), .O(n4664));
  orx   g04181(.a(n4664), .b(n4663), .O(n4665));
  orx   g04182(.a(n4665), .b(n4304), .O(n4666));
  invx  g04183(.a(n4666), .O(n4667));
  andx  g04184(.a(n4665), .b(n4304), .O(n4668));
  orx   g04185(.a(n4668), .b(n4667), .O(n4669));
  andx  g04186(.a(n3721), .b(n214), .O(n4670));
  orx   g04187(.a(n4670), .b(n4661), .O(n4671));
  andx  g04188(.a(n4671), .b(n4669), .O(n4672));
  orx   g04189(.a(n4672), .b(n4662), .O(n4673));
  andx  g04190(.a(n4673), .b(n4063), .O(n4674));
  andx  g04191(.a(n4436), .b(n4432), .O(n4675));
  andx  g04192(.a(n4435), .b(n4431), .O(n4676));
  orx   g04193(.a(n4676), .b(n4675), .O(n4677));
  andx  g04194(.a(n4677), .b(n4296), .O(n4678));
  invx  g04195(.a(n4678), .O(n4679));
  orx   g04196(.a(n4677), .b(n4296), .O(n4680));
  andx  g04197(.a(n4680), .b(n4679), .O(n4681));
  andx  g04198(.a(n4063), .b(n214), .O(n4682));
  orx   g04199(.a(n4682), .b(n4673), .O(n4683));
  andx  g04200(.a(n4683), .b(n4681), .O(n4684));
  orx   g04201(.a(n4684), .b(n4674), .O(n4685));
  andx  g04202(.a(n4685), .b(n4114), .O(n4686));
  andx  g04203(.a(n4449), .b(n4439), .O(n4687));
  andx  g04204(.a(n4448), .b(n4451), .O(n4688));
  orx   g04205(.a(n4688), .b(n4687), .O(n4689));
  invx  g04206(.a(n4689), .O(n4690));
  andx  g04207(.a(n4690), .b(n4446), .O(n4691));
  andx  g04208(.a(n4689), .b(n4452), .O(n4692));
  orx   g04209(.a(n4692), .b(n4691), .O(n4693));
  andx  g04210(.a(n4114), .b(n214), .O(n4694));
  orx   g04211(.a(n4694), .b(n4685), .O(n4695));
  andx  g04212(.a(n4695), .b(n4693), .O(n4696));
  orx   g04213(.a(n4696), .b(n4686), .O(n4697));
  andx  g04214(.a(n4697), .b(n4490), .O(n4698));
  andx  g04215(.a(n4461), .b(n4456), .O(n4699));
  andx  g04216(.a(n4460), .b(n4455), .O(n4700));
  orx   g04217(.a(n4700), .b(n4699), .O(n4701));
  andx  g04218(.a(n4701), .b(n4287), .O(n4702));
  invx  g04219(.a(n4702), .O(n4703));
  orx   g04220(.a(n4701), .b(n4287), .O(n4704));
  andx  g04221(.a(n4704), .b(n4703), .O(n4705));
  invx  g04222(.a(n4705), .O(n4706));
  andx  g04223(.a(n214), .b(n4706), .O(n4709));
  orx   g04224(.a(n4709), .b(n4698), .O(n4710));
  invx  g04225(.a(n4710), .O(n4716));
  andx  g04226(.a(n4716), .b(n4499), .O(n4717));
  invx  g04227(.a(n4499), .O(n4718));
  orx   g04228(.a(n4984), .b(n4717), .O(n4720));
  invx  g04229(.a(n4720), .O(n4721));
  invx  g04230(.a(n4698), .O(n4722));
  andx  g04231(.a(n214), .b(n4722), .O(n4723));
  invx  g04232(.a(n4723), .O(n4724));
  andx  g04233(.a(n4724), .b(n4705), .O(n4725));
  andx  g04234(.a(n4723), .b(n4706), .O(n4726));
  orx   g04235(.a(n4726), .b(n4725), .O(n4727));
  invx  g04236(.a(n4727), .O(n4728));
  invx  g04237(.a(n4693), .O(n4732));
  invx  g04238(.a(n4686), .O(n4733));
  andx  g04239(.a(n4695), .b(n4733), .O(n4734));
  invx  g04240(.a(n4734), .O(n4735));
  andx  g04241(.a(n4735), .b(n4732), .O(n4736));
  andx  g04242(.a(n4734), .b(n4693), .O(n4737));
  orx   g04243(.a(n4737), .b(n4736), .O(n4738));
  invx  g04244(.a(n4674), .O(n4739));
  andx  g04245(.a(n4683), .b(n4739), .O(n4740));
  orx   g04246(.a(n4740), .b(n4681), .O(n4741));
  andx  g04247(.a(n4740), .b(n4681), .O(n4742));
  invx  g04248(.a(n4742), .O(n4743));
  andx  g04249(.a(n4743), .b(n4741), .O(n4744));
  invx  g04250(.a(n4668), .O(n4745));
  andx  g04251(.a(n4745), .b(n4666), .O(n4746));
  invx  g04252(.a(n4662), .O(n4747));
  andx  g04253(.a(n4671), .b(n4747), .O(n4748));
  invx  g04254(.a(n4748), .O(n4749));
  andx  g04255(.a(n4749), .b(n4746), .O(n4750));
  andx  g04256(.a(n4748), .b(n4669), .O(n4751));
  orx   g04257(.a(n4751), .b(n4750), .O(n4752));
  andx  g04258(.a(n4659), .b(n4647), .O(n4753));
  orx   g04259(.a(n4753), .b(n4655), .O(n4754));
  invx  g04260(.a(n4655), .O(n4755));
  orx   g04261(.a(n4658), .b(n4648), .O(n4756));
  orx   g04262(.a(n4756), .b(n4755), .O(n4757));
  andx  g04263(.a(n4757), .b(n4754), .O(n4758));
  orx   g04264(.a(n4632), .b(n4627), .O(n4759));
  andx  g04265(.a(n4632), .b(n4627), .O(n4760));
  invx  g04266(.a(n4760), .O(n4761));
  andx  g04267(.a(n4761), .b(n4759), .O(n4762));
  orx   g04268(.a(n4762), .b(n4633), .O(n4763));
  invx  g04269(.a(n4759), .O(n4764));
  orx   g04270(.a(n4760), .b(n4764), .O(n4765));
  orx   g04271(.a(n4765), .b(n4547), .O(n4766));
  andx  g04272(.a(n4766), .b(n4763), .O(n4767));
  andx  g04273(.a(n4607), .b(n4603), .O(n4768));
  andx  g04274(.a(n4606), .b(n4608), .O(n4769));
  orx   g04275(.a(n4769), .b(n4768), .O(n4770));
  andx  g04276(.a(n4770), .b(n4573), .O(n4771));
  invx  g04277(.a(n4771), .O(n4772));
  orx   g04278(.a(n4770), .b(n4573), .O(n4773));
  andx  g04279(.a(n4773), .b(n4772), .O(n4774));
  invx  g04280(.a(n4588), .O(n4775));
  andx  g04281(.a(n4601), .b(n4775), .O(n4776));
  invx  g04282(.a(n4776), .O(n4777));
  andx  g04283(.a(n4777), .b(n4599), .O(n4778));
  invx  g04284(.a(n4599), .O(n4779));
  andx  g04285(.a(n4776), .b(n4779), .O(n4780));
  orx   g04286(.a(n4780), .b(n4778), .O(n4781));
  andx  g04287(.a(n3230), .b(n250), .O(n4782));
  invx  g04288(.a(n4582), .O(n4783));
  andx  g04289(.a(n4783), .b(n4581), .O(n4784));
  invx  g04290(.a(n4581), .O(n4785));
  andx  g04291(.a(n4582), .b(n4785), .O(n4786));
  orx   g04292(.a(n4786), .b(n4784), .O(n4787));
  andx  g04293(.a(n4787), .b(n4782), .O(n4788));
  andx  g04294(.a(n1790), .b(n214), .O(n4789));
  andx  g04295(.a(n3258), .b(n250), .O(n4790));
  andx  g04296(.a(n4790), .b(n4789), .O(n4791));
  andx  g04297(.a(n4791), .b(n4782), .O(n4792));
  andx  g04298(.a(n4791), .b(n4787), .O(n4793));
  orx   g04299(.a(n4793), .b(n4792), .O(n4794));
  orx   g04300(.a(n4794), .b(n4788), .O(n4795));
  andx  g04301(.a(n4795), .b(n3221), .O(n4796));
  invx  g04302(.a(n4583), .O(n4797));
  andx  g04303(.a(n4797), .b(n4574), .O(n4798));
  invx  g04304(.a(n4798), .O(n4799));
  orx   g04305(.a(n4797), .b(n4574), .O(n4800));
  andx  g04306(.a(n4800), .b(n4799), .O(n4801));
  andx  g04307(.a(n4575), .b(n4577), .O(n4802));
  orx   g04308(.a(n4802), .b(n4337), .O(n4803));
  andx  g04309(.a(n4803), .b(n4801), .O(n4804));
  invx  g04310(.a(n4804), .O(n4805));
  orx   g04311(.a(n4803), .b(n4801), .O(n4806));
  andx  g04312(.a(n4806), .b(n4805), .O(n4807));
  andx  g04313(.a(n3221), .b(n250), .O(n4808));
  orx   g04314(.a(n4808), .b(n4795), .O(n4809));
  andx  g04315(.a(n4809), .b(n4807), .O(n4810));
  orx   g04316(.a(n4810), .b(n4796), .O(n4811));
  andx  g04317(.a(n4811), .b(n4781), .O(n4812));
  andx  g04318(.a(n3210), .b(n250), .O(n4813));
  orx   g04319(.a(n4811), .b(n4781), .O(n4814));
  andx  g04320(.a(n4814), .b(n4813), .O(n4815));
  orx   g04321(.a(n4815), .b(n4812), .O(n4816));
  andx  g04322(.a(n4816), .b(n4774), .O(n4817));
  invx  g04323(.a(n4817), .O(n4818));
  invx  g04324(.a(n4773), .O(n4819));
  orx   g04325(.a(n4819), .b(n4771), .O(n4820));
  invx  g04326(.a(n4812), .O(n4821));
  invx  g04327(.a(n4813), .O(n4822));
  orx   g04328(.a(n4776), .b(n4779), .O(n4823));
  orx   g04329(.a(n4777), .b(n4599), .O(n4824));
  andx  g04330(.a(n4824), .b(n4823), .O(n4825));
  invx  g04331(.a(n4811), .O(n4826));
  andx  g04332(.a(n4826), .b(n4825), .O(n4827));
  orx   g04333(.a(n4827), .b(n4822), .O(n4828));
  andx  g04334(.a(n4828), .b(n4821), .O(n4829));
  andx  g04335(.a(n4829), .b(n4820), .O(n4830));
  andx  g04336(.a(n3284), .b(n250), .O(n4831));
  invx  g04337(.a(n4831), .O(n4832));
  orx   g04338(.a(n4832), .b(n4830), .O(n4833));
  andx  g04339(.a(n4833), .b(n4818), .O(n4834));
  orx   g04340(.a(n4616), .b(n4611), .O(n4835));
  andx  g04341(.a(n4616), .b(n4611), .O(n4836));
  invx  g04342(.a(n4836), .O(n4837));
  andx  g04343(.a(n4837), .b(n4835), .O(n4838));
  orx   g04344(.a(n4838), .b(n4565), .O(n4839));
  invx  g04345(.a(n4835), .O(n4840));
  orx   g04346(.a(n4836), .b(n4840), .O(n4841));
  orx   g04347(.a(n4841), .b(n4564), .O(n4842));
  andx  g04348(.a(n4842), .b(n4839), .O(n4843));
  andx  g04349(.a(n4843), .b(n4834), .O(n4844));
  andx  g04350(.a(n3180), .b(n250), .O(n4845));
  invx  g04351(.a(n4845), .O(n4846));
  orx   g04352(.a(n4846), .b(n4844), .O(n4847));
  orx   g04353(.a(n4816), .b(n4774), .O(n4848));
  andx  g04354(.a(n4831), .b(n4848), .O(n4849));
  orx   g04355(.a(n4849), .b(n4817), .O(n4850));
  andx  g04356(.a(n4841), .b(n4564), .O(n4851));
  andx  g04357(.a(n4838), .b(n4565), .O(n4852));
  orx   g04358(.a(n4852), .b(n4851), .O(n4853));
  andx  g04359(.a(n4853), .b(n4850), .O(n4854));
  invx  g04360(.a(n4854), .O(n4855));
  andx  g04361(.a(n4855), .b(n4847), .O(n4856));
  andx  g04362(.a(n4624), .b(n4619), .O(n4857));
  orx   g04363(.a(n4624), .b(n4619), .O(n4858));
  invx  g04364(.a(n4858), .O(n4859));
  orx   g04365(.a(n4859), .b(n4857), .O(n4860));
  andx  g04366(.a(n4860), .b(n4555), .O(n4861));
  invx  g04367(.a(n4857), .O(n4862));
  andx  g04368(.a(n4858), .b(n4862), .O(n4863));
  andx  g04369(.a(n4863), .b(n4556), .O(n4864));
  orx   g04370(.a(n4864), .b(n4861), .O(n4865));
  andx  g04371(.a(n4865), .b(n4856), .O(n4866));
  andx  g04372(.a(n3429), .b(n250), .O(n4867));
  invx  g04373(.a(n4867), .O(n4868));
  andx  g04374(.a(n4868), .b(n4856), .O(n4869));
  andx  g04375(.a(n4868), .b(n4865), .O(n4870));
  orx   g04376(.a(n4870), .b(n4869), .O(n4871));
  orx   g04377(.a(n4871), .b(n4866), .O(n4872));
  andx  g04378(.a(n4872), .b(n4767), .O(n4873));
  andx  g04379(.a(n3171), .b(n250), .O(n4874));
  invx  g04380(.a(n4874), .O(n4875));
  andx  g04381(.a(n4875), .b(n4767), .O(n4876));
  andx  g04382(.a(n4875), .b(n4872), .O(n4877));
  orx   g04383(.a(n4877), .b(n4876), .O(n4878));
  orx   g04384(.a(n4878), .b(n4873), .O(n4879));
  orx   g04385(.a(n4636), .b(n4532), .O(n4880));
  andx  g04386(.a(n4636), .b(n4532), .O(n4881));
  invx  g04387(.a(n4881), .O(n4882));
  andx  g04388(.a(n4882), .b(n4880), .O(n4883));
  andx  g04389(.a(n4883), .b(n4528), .O(n4884));
  invx  g04390(.a(n4880), .O(n4885));
  orx   g04391(.a(n4881), .b(n4885), .O(n4886));
  andx  g04392(.a(n4886), .b(n4527), .O(n4887));
  orx   g04393(.a(n4887), .b(n4884), .O(n4888));
  andx  g04394(.a(n4888), .b(n4879), .O(n4889));
  andx  g04395(.a(n3413), .b(n250), .O(n4890));
  invx  g04396(.a(n4890), .O(n4891));
  orx   g04397(.a(n4891), .b(n4889), .O(n4892));
  invx  g04398(.a(n4873), .O(n4893));
  andx  g04399(.a(n4765), .b(n4547), .O(n4894));
  andx  g04400(.a(n4762), .b(n4633), .O(n4895));
  orx   g04401(.a(n4895), .b(n4894), .O(n4896));
  orx   g04402(.a(n4874), .b(n4896), .O(n4897));
  invx  g04403(.a(n4877), .O(n4898));
  andx  g04404(.a(n4898), .b(n4897), .O(n4899));
  andx  g04405(.a(n4899), .b(n4893), .O(n4900));
  orx   g04406(.a(n4886), .b(n4527), .O(n4901));
  orx   g04407(.a(n4883), .b(n4528), .O(n4902));
  andx  g04408(.a(n4902), .b(n4901), .O(n4903));
  andx  g04409(.a(n4903), .b(n4900), .O(n4904));
  invx  g04410(.a(n4904), .O(n4905));
  andx  g04411(.a(n4905), .b(n4892), .O(n4906));
  orx   g04412(.a(n4643), .b(n4638), .O(n4907));
  andx  g04413(.a(n4643), .b(n4638), .O(n4908));
  invx  g04414(.a(n4908), .O(n4909));
  andx  g04415(.a(n4909), .b(n4907), .O(n4910));
  orx   g04416(.a(n4910), .b(n4517), .O(n4911));
  invx  g04417(.a(n4907), .O(n4912));
  orx   g04418(.a(n4908), .b(n4912), .O(n4913));
  orx   g04419(.a(n4913), .b(n4518), .O(n4914));
  andx  g04420(.a(n4914), .b(n4911), .O(n4915));
  andx  g04421(.a(n4915), .b(n4906), .O(n4916));
  invx  g04422(.a(n4916), .O(n4917));
  orx   g04423(.a(n4903), .b(n4900), .O(n4918));
  andx  g04424(.a(n4890), .b(n4918), .O(n4919));
  orx   g04425(.a(n4904), .b(n4919), .O(n4920));
  andx  g04426(.a(n3645), .b(n250), .O(n4921));
  orx   g04427(.a(n4921), .b(n4920), .O(n4922));
  andx  g04428(.a(n4913), .b(n4518), .O(n4923));
  andx  g04429(.a(n4910), .b(n4517), .O(n4924));
  orx   g04430(.a(n4924), .b(n4923), .O(n4925));
  orx   g04431(.a(n4921), .b(n4925), .O(n4926));
  andx  g04432(.a(n4926), .b(n4922), .O(n4927));
  andx  g04433(.a(n4927), .b(n4917), .O(n4928));
  andx  g04434(.a(n4928), .b(n4758), .O(n4929));
  invx  g04435(.a(n4929), .O(n4930));
  andx  g04436(.a(n3721), .b(n250), .O(n4931));
  invx  g04437(.a(n4931), .O(n4932));
  andx  g04438(.a(n4756), .b(n4755), .O(n4933));
  andx  g04439(.a(n4753), .b(n4655), .O(n4934));
  orx   g04440(.a(n4934), .b(n4933), .O(n4935));
  invx  g04441(.a(n4921), .O(n4936));
  andx  g04442(.a(n4936), .b(n4906), .O(n4937));
  andx  g04443(.a(n4936), .b(n4915), .O(n4938));
  orx   g04444(.a(n4938), .b(n4937), .O(n4939));
  orx   g04445(.a(n4939), .b(n4916), .O(n4940));
  andx  g04446(.a(n4940), .b(n4935), .O(n4941));
  orx   g04447(.a(n4941), .b(n4932), .O(n4942));
  andx  g04448(.a(n4942), .b(n4930), .O(n4943));
  andx  g04449(.a(n4943), .b(n4752), .O(n4944));
  andx  g04450(.a(n4063), .b(n250), .O(n4945));
  invx  g04451(.a(n4945), .O(n4946));
  orx   g04452(.a(n4946), .b(n4944), .O(n4947));
  orx   g04453(.a(n4748), .b(n4669), .O(n4948));
  orx   g04454(.a(n4749), .b(n4746), .O(n4949));
  andx  g04455(.a(n4949), .b(n4948), .O(n4950));
  orx   g04456(.a(n4928), .b(n4758), .O(n4951));
  andx  g04457(.a(n4951), .b(n4931), .O(n4952));
  orx   g04458(.a(n4952), .b(n4929), .O(n4953));
  andx  g04459(.a(n4953), .b(n4950), .O(n4954));
  invx  g04460(.a(n4954), .O(n4955));
  andx  g04461(.a(n4955), .b(n4947), .O(n4956));
  invx  g04462(.a(n4956), .O(n4957));
  andx  g04463(.a(n4957), .b(n4744), .O(n4958));
  invx  g04464(.a(n4958), .O(n4959));
  invx  g04465(.a(n4741), .O(n4960));
  orx   g04466(.a(n4742), .b(n4960), .O(n4961));
  andx  g04467(.a(n4956), .b(n4961), .O(n4962));
  andx  g04468(.a(n4114), .b(n250), .O(n4963));
  invx  g04469(.a(n4963), .O(n4964));
  orx   g04470(.a(n4964), .b(n4962), .O(n4965));
  andx  g04471(.a(n4965), .b(n4959), .O(n4966));
  andx  g04472(.a(n4966), .b(n4738), .O(n4967));
  andx  g04473(.a(n4490), .b(n250), .O(n4968));
  invx  g04474(.a(n4968), .O(n4969));
  orx   g04475(.a(n4969), .b(n4967), .O(n4970));
  invx  g04476(.a(n4738), .O(n4971));
  orx   g04477(.a(n4957), .b(n4744), .O(n4972));
  andx  g04478(.a(n4963), .b(n4972), .O(n4973));
  orx   g04479(.a(n4973), .b(n4958), .O(n4974));
  andx  g04480(.a(n4974), .b(n4971), .O(n4975));
  invx  g04481(.a(n4975), .O(n4976));
  andx  g04482(.a(n4976), .b(n4970), .O(n4977));
  orx   g04483(.a(n4727), .b(n4977), .O(n4980));
  andx  g04484(.a(n5391), .b(n4721), .O(n4983));
  andx  g04485(.a(n4710), .b(n4718), .O(n4984));
  invx  g04486(.a(n4984), .O(n4986));
  andx  g04487(.a(n3403), .b(n3313), .O(n4987));
  andx  g04488(.a(n4987), .b(n3158), .O(n4988));
  orx   g04489(.a(n4988), .b(n3562), .O(n4989));
  andx  g04490(.a(n3645), .b(n827), .O(n4990));
  orx   g04491(.a(n4990), .b(n4989), .O(n4991));
  andx  g04492(.a(n4989), .b(n827), .O(n4992));
  andx  g04493(.a(n4992), .b(n3645), .O(n4993));
  invx  g04494(.a(n4993), .O(n4994));
  andx  g04495(.a(n4994), .b(n4991), .O(n4995));
  invx  g04496(.a(n4995), .O(n4996));
  andx  g04497(.a(n3311), .b(n3171), .O(n4997));
  invx  g04498(.a(n4997), .O(n4998));
  andx  g04499(.a(n3310), .b(n3307), .O(n4999));
  orx   g04500(.a(n4999), .b(n4989), .O(n5000));
  andx  g04501(.a(n5000), .b(n4998), .O(n5001));
  invx  g04502(.a(n5001), .O(n5002));
  andx  g04503(.a(n5002), .b(n4996), .O(n5003));
  andx  g04504(.a(n5001), .b(n4995), .O(n5004));
  orx   g04505(.a(n5004), .b(n5003), .O(n5005));
  andx  g04506(.a(n3649), .b(n3424), .O(n5006));
  invx  g04507(.a(n5006), .O(n5007));
  andx  g04508(.a(n3559), .b(n3425), .O(n5008));
  orx   g04509(.a(n5008), .b(n3647), .O(n5009));
  andx  g04510(.a(n5009), .b(n5007), .O(n5010));
  invx  g04511(.a(n5010), .O(n5011));
  andx  g04512(.a(n3721), .b(n299), .O(n5012));
  invx  g04513(.a(n5012), .O(n5013));
  andx  g04514(.a(n5013), .b(n5011), .O(n5014));
  andx  g04515(.a(n5012), .b(n5010), .O(n5015));
  orx   g04516(.a(n5015), .b(n5014), .O(n5016));
  andx  g04517(.a(n5016), .b(n5005), .O(n5017));
  invx  g04518(.a(n5017), .O(n5018));
  orx   g04519(.a(n5016), .b(n5005), .O(n5019));
  andx  g04520(.a(n5019), .b(n5018), .O(n5020));
  andx  g04521(.a(n3847), .b(n3655), .O(n5021));
  orx   g04522(.a(n5021), .b(n3844), .O(n5022));
  andx  g04523(.a(n5022), .b(n4063), .O(n5023));
  invx  g04524(.a(n5023), .O(n5024));
  andx  g04525(.a(n4063), .b(n338), .O(n5025));
  orx   g04526(.a(n5025), .b(n5022), .O(n5026));
  andx  g04527(.a(n5026), .b(n5024), .O(n5027));
  invx  g04528(.a(n5027), .O(n5028));
  andx  g04529(.a(n5028), .b(n5020), .O(n5029));
  invx  g04530(.a(n5020), .O(n5030));
  andx  g04531(.a(n5027), .b(n5030), .O(n5031));
  orx   g04532(.a(n5031), .b(n5029), .O(n5032));
  andx  g04533(.a(n4014), .b(n3852), .O(n5033));
  orx   g04534(.a(n5033), .b(n4065), .O(n5034));
  orx   g04535(.a(n4014), .b(n3852), .O(n5035));
  andx  g04536(.a(n5035), .b(n5034), .O(n5036));
  invx  g04537(.a(n5036), .O(n5037));
  andx  g04538(.a(n4114), .b(n376), .O(n5038));
  invx  g04539(.a(n5038), .O(n5039));
  andx  g04540(.a(n5039), .b(n5037), .O(n5040));
  andx  g04541(.a(n5038), .b(n5036), .O(n5041));
  orx   g04542(.a(n5041), .b(n5040), .O(n5042));
  andx  g04543(.a(n5042), .b(n5032), .O(n5043));
  invx  g04544(.a(n5043), .O(n5044));
  orx   g04545(.a(n5042), .b(n5032), .O(n5045));
  andx  g04546(.a(n5045), .b(n5044), .O(n5046));
  andx  g04547(.a(n4275), .b(n4279), .O(n5047));
  orx   g04548(.a(n5047), .b(n4272), .O(n5048));
  andx  g04549(.a(n5048), .b(n4490), .O(n5049));
  invx  g04550(.a(n5049), .O(n5050));
  andx  g04551(.a(n4490), .b(n438), .O(n5051));
  orx   g04552(.a(n5051), .b(n5048), .O(n5052));
  andx  g04553(.a(n5052), .b(n5050), .O(n5053));
  invx  g04554(.a(n5053), .O(n5054));
  andx  g04555(.a(n5054), .b(n5046), .O(n5055));
  invx  g04556(.a(n5046), .O(n5056));
  andx  g04557(.a(n5053), .b(n5056), .O(n5057));
  orx   g04558(.a(n5057), .b(n5055), .O(n5058));
  andx  g04559(.a(n2724), .b(n252), .O(n5059));
  invx  g04560(.a(n5059), .O(n5060));
  andx  g04561(.a(n4463), .b(n4281), .O(n5061));
  orx   g04562(.a(n5061), .b(n4492), .O(n5062));
  orx   g04563(.a(n4463), .b(n4281), .O(n5063));
  andx  g04564(.a(n5063), .b(n5062), .O(n5064));
  invx  g04565(.a(n5064), .O(n5065));
  andx  g04566(.a(n5065), .b(n5060), .O(n5066));
  andx  g04567(.a(n5066), .b(n5058), .O(n5069));
  invx  g04568(.a(n5069), .O(n5070));
  orx   g04569(.a(n5066), .b(n5058), .O(n5071));
  andx  g04570(.a(n5071), .b(n5070), .O(n5072));
  invx  g04571(.a(n5072), .O(n5073));
  andx  g04572(.a(n5073), .b(n4986), .O(n5074));
  andx  g04573(.a(n5072), .b(n4984), .O(n5075));
  orx   g04574(.a(n5075), .b(n5074), .O(n5076));
  andx  g04575(.a(n5076), .b(n4983), .O(n5077));
  andx  g04576(.a(n5073), .b(n4984), .O(n5078));
  orx   g04577(.a(n5078), .b(n5077), .O(n5079));
  orx   g04578(.a(n4977), .b(n3011), .O(n5080));
  invx  g04579(.a(n5080), .O(n5081));
  andx  g04580(.a(n4977), .b(n3011), .O(n5082));
  orx   g04581(.a(n5082), .b(n5081), .O(n5083));
  invx  g04582(.a(n5082), .O(n5085));
  andx  g04583(.a(n5085), .b(n5080), .O(n5086));
  orx   g04584(.a(n5086), .b(n4728), .O(n5087));
  andx  g04585(.a(n5087), .b(n4980), .O(n5088));
  andx  g04586(.a(n4921), .b(n4920), .O(n5098));
  orx   g04587(.a(n5098), .b(n4937), .O(n5099));
  orx   g04588(.a(n5099), .b(n4915), .O(n5100));
  orx   g04589(.a(n4936), .b(n4906), .O(n5104));
  andx  g04590(.a(n5104), .b(n4922), .O(n5105));
  orx   g04591(.a(n5105), .b(n4925), .O(n5106));
  andx  g04592(.a(n5106), .b(n5100), .O(n5107));
  andx  g04593(.a(n4874), .b(n4872), .O(n5108));
  invx  g04594(.a(n4866), .O(n5109));
  orx   g04595(.a(n4853), .b(n4850), .O(n5110));
  andx  g04596(.a(n4845), .b(n5110), .O(n5111));
  orx   g04597(.a(n4854), .b(n5111), .O(n5112));
  orx   g04598(.a(n4867), .b(n5112), .O(n5113));
  orx   g04599(.a(n4863), .b(n4556), .O(n5114));
  orx   g04600(.a(n4860), .b(n4555), .O(n5115));
  andx  g04601(.a(n5115), .b(n5114), .O(n5116));
  orx   g04602(.a(n4867), .b(n5116), .O(n5117));
  andx  g04603(.a(n5117), .b(n5113), .O(n5118));
  andx  g04604(.a(n5118), .b(n5109), .O(n5119));
  andx  g04605(.a(n4875), .b(n5119), .O(n5120));
  orx   g04606(.a(n5120), .b(n5108), .O(n5121));
  andx  g04607(.a(n4896), .b(n5121), .O(n5131));
  orx   g04608(.a(n4875), .b(n5119), .O(n5132));
  orx   g04609(.a(n4874), .b(n4872), .O(n5133));
  andx  g04610(.a(n5133), .b(n5132), .O(n5134));
  andx  g04611(.a(n4767), .b(n5134), .O(n5138));
  orx   g04612(.a(n5138), .b(n5131), .O(n5139));
  andx  g04613(.a(n4867), .b(n5112), .O(n5143));
  orx   g04614(.a(n5143), .b(n4869), .O(n5144));
  orx   g04615(.a(n5144), .b(n4865), .O(n5145));
  orx   g04616(.a(n4868), .b(n4856), .O(n5149));
  andx  g04617(.a(n5149), .b(n5113), .O(n5150));
  orx   g04618(.a(n5150), .b(n5116), .O(n5151));
  andx  g04619(.a(n5151), .b(n5145), .O(n5152));
  orx   g04620(.a(n4831), .b(n4829), .O(n5153));
  orx   g04621(.a(n4832), .b(n4816), .O(n5154));
  andx  g04622(.a(n5154), .b(n5153), .O(n5155));
  orx   g04623(.a(n5155), .b(n4774), .O(n5156));
  andx  g04624(.a(n4832), .b(n4816), .O(n5157));
  andx  g04625(.a(n4831), .b(n4829), .O(n5158));
  orx   g04626(.a(n5158), .b(n5157), .O(n5159));
  orx   g04627(.a(n5159), .b(n4820), .O(n5160));
  andx  g04628(.a(n5160), .b(n5156), .O(n5161));
  andx  g04629(.a(n4822), .b(n4811), .O(n5162));
  invx  g04630(.a(n5162), .O(n5163));
  orx   g04631(.a(n4822), .b(n4811), .O(n5164));
  andx  g04632(.a(n5164), .b(n5163), .O(n5165));
  orx   g04633(.a(n5165), .b(n4825), .O(n5166));
  invx  g04634(.a(n5164), .O(n5167));
  orx   g04635(.a(n5167), .b(n5162), .O(n5168));
  orx   g04636(.a(n5168), .b(n4781), .O(n5169));
  andx  g04637(.a(n5169), .b(n5166), .O(n5170));
  invx  g04638(.a(n4809), .O(n5171));
  orx   g04639(.a(n5171), .b(n4796), .O(n5172));
  andx  g04640(.a(n5172), .b(n4807), .O(n5173));
  invx  g04641(.a(n4806), .O(n5174));
  orx   g04642(.a(n5174), .b(n4804), .O(n5175));
  invx  g04643(.a(n4796), .O(n5176));
  andx  g04644(.a(n4809), .b(n5176), .O(n5177));
  andx  g04645(.a(n5177), .b(n5175), .O(n5178));
  orx   g04646(.a(n5178), .b(n5173), .O(n5179));
  andx  g04647(.a(n3230), .b(n403), .O(n5180));
  orx   g04648(.a(n3490), .b(n179), .O(n5181));
  andx  g04649(.a(n5181), .b(n4789), .O(n5182));
  invx  g04650(.a(n4789), .O(n5183));
  andx  g04651(.a(n4790), .b(n5183), .O(n5184));
  orx   g04652(.a(n5184), .b(n5182), .O(n5185));
  andx  g04653(.a(n5185), .b(n5180), .O(n5186));
  andx  g04654(.a(n3258), .b(n403), .O(n5187));
  andx  g04655(.a(n1790), .b(n250), .O(n5188));
  andx  g04656(.a(n5188), .b(n5187), .O(n5189));
  andx  g04657(.a(n5189), .b(n5180), .O(n5190));
  andx  g04658(.a(n5189), .b(n5185), .O(n5191));
  orx   g04659(.a(n5191), .b(n5190), .O(n5192));
  orx   g04660(.a(n5192), .b(n5186), .O(n5193));
  andx  g04661(.a(n5193), .b(n3221), .O(n5194));
  invx  g04662(.a(n4791), .O(n5195));
  andx  g04663(.a(n5195), .b(n4782), .O(n5196));
  orx   g04664(.a(n3239), .b(n179), .O(n5197));
  andx  g04665(.a(n4791), .b(n5197), .O(n5198));
  orx   g04666(.a(n5198), .b(n5196), .O(n5199));
  andx  g04667(.a(n4783), .b(n4785), .O(n5200));
  orx   g04668(.a(n5200), .b(n4583), .O(n5201));
  orx   g04669(.a(n4787), .b(n5199), .O(n5203));
  orx   g04670(.a(n4791), .b(n5197), .O(n5204));
  orx   g04671(.a(n5195), .b(n4782), .O(n5205));
  andx  g04672(.a(n5205), .b(n5204), .O(n5206));
  orx   g04673(.a(n5201), .b(n5206), .O(n5207));
  andx  g04674(.a(n5207), .b(n5203), .O(n5208));
  andx  g04675(.a(n3221), .b(n403), .O(n5209));
  orx   g04676(.a(n5209), .b(n5193), .O(n5210));
  andx  g04677(.a(n5210), .b(n5208), .O(n5211));
  orx   g04678(.a(n5211), .b(n5194), .O(n5212));
  andx  g04679(.a(n5212), .b(n5179), .O(n5213));
  andx  g04680(.a(n3210), .b(n403), .O(n5214));
  orx   g04681(.a(n5212), .b(n5179), .O(n5215));
  andx  g04682(.a(n5215), .b(n5214), .O(n5216));
  orx   g04683(.a(n5216), .b(n5213), .O(n5217));
  andx  g04684(.a(n5217), .b(n5170), .O(n5218));
  invx  g04685(.a(n5218), .O(n5219));
  andx  g04686(.a(n5168), .b(n4781), .O(n5220));
  andx  g04687(.a(n5165), .b(n4825), .O(n5221));
  orx   g04688(.a(n5221), .b(n5220), .O(n5222));
  invx  g04689(.a(n5213), .O(n5223));
  invx  g04690(.a(n5214), .O(n5224));
  orx   g04691(.a(n5177), .b(n5175), .O(n5225));
  orx   g04692(.a(n5172), .b(n4807), .O(n5226));
  andx  g04693(.a(n5226), .b(n5225), .O(n5227));
  invx  g04694(.a(n5212), .O(n5228));
  andx  g04695(.a(n5228), .b(n5227), .O(n5229));
  orx   g04696(.a(n5229), .b(n5224), .O(n5230));
  andx  g04697(.a(n5230), .b(n5223), .O(n5231));
  andx  g04698(.a(n5231), .b(n5222), .O(n5232));
  andx  g04699(.a(n3284), .b(n403), .O(n5233));
  invx  g04700(.a(n5233), .O(n5234));
  orx   g04701(.a(n5234), .b(n5232), .O(n5235));
  andx  g04702(.a(n5235), .b(n5219), .O(n5236));
  andx  g04703(.a(n5236), .b(n5161), .O(n5237));
  andx  g04704(.a(n3180), .b(n403), .O(n5238));
  invx  g04705(.a(n5238), .O(n5239));
  orx   g04706(.a(n5239), .b(n5237), .O(n5240));
  andx  g04707(.a(n5159), .b(n4820), .O(n5241));
  andx  g04708(.a(n5155), .b(n4774), .O(n5242));
  orx   g04709(.a(n5242), .b(n5241), .O(n5243));
  orx   g04710(.a(n5217), .b(n5170), .O(n5244));
  andx  g04711(.a(n5233), .b(n5244), .O(n5245));
  orx   g04712(.a(n5245), .b(n5218), .O(n5246));
  andx  g04713(.a(n5246), .b(n5243), .O(n5247));
  invx  g04714(.a(n5247), .O(n5248));
  andx  g04715(.a(n5248), .b(n5240), .O(n5249));
  andx  g04716(.a(n4846), .b(n4834), .O(n5250));
  andx  g04717(.a(n4845), .b(n4850), .O(n5251));
  orx   g04718(.a(n5251), .b(n5250), .O(n5252));
  andx  g04719(.a(n5252), .b(n4843), .O(n5253));
  orx   g04720(.a(n4845), .b(n4850), .O(n5254));
  orx   g04721(.a(n4846), .b(n4834), .O(n5255));
  andx  g04722(.a(n5255), .b(n5254), .O(n5256));
  andx  g04723(.a(n5256), .b(n4853), .O(n5257));
  orx   g04724(.a(n5257), .b(n5253), .O(n5258));
  andx  g04725(.a(n5258), .b(n5249), .O(n5259));
  invx  g04726(.a(n5259), .O(n5260));
  orx   g04727(.a(n5246), .b(n5243), .O(n5261));
  andx  g04728(.a(n5238), .b(n5261), .O(n5262));
  orx   g04729(.a(n5247), .b(n5262), .O(n5263));
  andx  g04730(.a(n3429), .b(n403), .O(n5264));
  orx   g04731(.a(n5264), .b(n5263), .O(n5265));
  orx   g04732(.a(n5256), .b(n4853), .O(n5266));
  orx   g04733(.a(n5252), .b(n4843), .O(n5267));
  andx  g04734(.a(n5267), .b(n5266), .O(n5268));
  orx   g04735(.a(n5264), .b(n5268), .O(n5269));
  andx  g04736(.a(n5269), .b(n5265), .O(n5270));
  andx  g04737(.a(n5270), .b(n5260), .O(n5271));
  andx  g04738(.a(n5271), .b(n5152), .O(n5272));
  invx  g04739(.a(n5272), .O(n5273));
  andx  g04740(.a(n3171), .b(n403), .O(n5274));
  invx  g04741(.a(n5274), .O(n5275));
  andx  g04742(.a(n5150), .b(n5116), .O(n5276));
  andx  g04743(.a(n5144), .b(n4865), .O(n5277));
  orx   g04744(.a(n5277), .b(n5276), .O(n5278));
  invx  g04745(.a(n5264), .O(n5279));
  andx  g04746(.a(n5279), .b(n5249), .O(n5280));
  andx  g04747(.a(n5279), .b(n5258), .O(n5281));
  orx   g04748(.a(n5281), .b(n5280), .O(n5282));
  orx   g04749(.a(n5282), .b(n5259), .O(n5283));
  andx  g04750(.a(n5283), .b(n5278), .O(n5284));
  orx   g04751(.a(n5284), .b(n5275), .O(n5285));
  andx  g04752(.a(n5285), .b(n5273), .O(n5286));
  andx  g04753(.a(n5286), .b(n5139), .O(n5287));
  andx  g04754(.a(n3413), .b(n403), .O(n5288));
  invx  g04755(.a(n5288), .O(n5289));
  orx   g04756(.a(n5289), .b(n5287), .O(n5290));
  orx   g04757(.a(n4767), .b(n5134), .O(n5291));
  orx   g04758(.a(n4896), .b(n5121), .O(n5292));
  andx  g04759(.a(n5292), .b(n5291), .O(n5293));
  orx   g04760(.a(n5271), .b(n5152), .O(n5294));
  andx  g04761(.a(n5294), .b(n5274), .O(n5295));
  orx   g04762(.a(n5295), .b(n5272), .O(n5296));
  andx  g04763(.a(n5296), .b(n5293), .O(n5297));
  invx  g04764(.a(n5297), .O(n5298));
  andx  g04765(.a(n5298), .b(n5290), .O(n5299));
  orx   g04766(.a(n4890), .b(n4879), .O(n5300));
  orx   g04767(.a(n4891), .b(n4900), .O(n5301));
  andx  g04768(.a(n5301), .b(n5300), .O(n5302));
  andx  g04769(.a(n5302), .b(n4888), .O(n5303));
  andx  g04770(.a(n4891), .b(n4900), .O(n5304));
  andx  g04771(.a(n4890), .b(n4879), .O(n5305));
  orx   g04772(.a(n5305), .b(n5304), .O(n5306));
  andx  g04773(.a(n5306), .b(n4903), .O(n5307));
  orx   g04774(.a(n5307), .b(n5303), .O(n5308));
  andx  g04775(.a(n5308), .b(n5299), .O(n5309));
  invx  g04776(.a(n5309), .O(n5310));
  orx   g04777(.a(n5296), .b(n5293), .O(n5311));
  andx  g04778(.a(n5288), .b(n5311), .O(n5312));
  orx   g04779(.a(n5297), .b(n5312), .O(n5313));
  andx  g04780(.a(n3645), .b(n403), .O(n5314));
  orx   g04781(.a(n5314), .b(n5313), .O(n5315));
  orx   g04782(.a(n5306), .b(n4903), .O(n5316));
  orx   g04783(.a(n5302), .b(n4888), .O(n5317));
  andx  g04784(.a(n5317), .b(n5316), .O(n5318));
  orx   g04785(.a(n5314), .b(n5318), .O(n5319));
  andx  g04786(.a(n5319), .b(n5315), .O(n5320));
  andx  g04787(.a(n5320), .b(n5310), .O(n5321));
  andx  g04788(.a(n5321), .b(n5107), .O(n5322));
  andx  g04789(.a(n3721), .b(n403), .O(n5323));
  orx   g04790(.a(n5321), .b(n5107), .O(n5324));
  andx  g04791(.a(n5324), .b(n5323), .O(n5325));
  orx   g04792(.a(n5325), .b(n5322), .O(n5326));
  andx  g04793(.a(n5326), .b(n4063), .O(n5327));
  orx   g04794(.a(n4932), .b(n4940), .O(n5328));
  orx   g04795(.a(n4931), .b(n4928), .O(n5329));
  andx  g04796(.a(n5329), .b(n5328), .O(n5330));
  andx  g04797(.a(n5330), .b(n4935), .O(n5331));
  andx  g04798(.a(n4931), .b(n4928), .O(n5332));
  andx  g04799(.a(n4932), .b(n4940), .O(n5333));
  orx   g04800(.a(n5333), .b(n5332), .O(n5334));
  andx  g04801(.a(n5334), .b(n4758), .O(n5335));
  orx   g04802(.a(n5335), .b(n5331), .O(n5336));
  andx  g04803(.a(n4063), .b(n403), .O(n5337));
  orx   g04804(.a(n5337), .b(n5326), .O(n5338));
  andx  g04805(.a(n5338), .b(n5336), .O(n5339));
  orx   g04806(.a(n5339), .b(n5327), .O(n5340));
  andx  g04807(.a(n5340), .b(n4114), .O(n5341));
  orx   g04808(.a(n4945), .b(n4953), .O(n5342));
  orx   g04809(.a(n4946), .b(n4943), .O(n5343));
  andx  g04810(.a(n5343), .b(n5342), .O(n5344));
  andx  g04811(.a(n5344), .b(n4752), .O(n5345));
  andx  g04812(.a(n4946), .b(n4943), .O(n5346));
  andx  g04813(.a(n4945), .b(n4953), .O(n5347));
  orx   g04814(.a(n5347), .b(n5346), .O(n5348));
  andx  g04815(.a(n5348), .b(n4950), .O(n5349));
  orx   g04816(.a(n5349), .b(n5345), .O(n5350));
  andx  g04817(.a(n4114), .b(n403), .O(n5351));
  orx   g04818(.a(n5351), .b(n5340), .O(n5352));
  andx  g04819(.a(n5352), .b(n5350), .O(n5353));
  orx   g04820(.a(n5353), .b(n5341), .O(n5354));
  andx  g04821(.a(n5354), .b(n4490), .O(n5355));
  orx   g04822(.a(n4963), .b(n4956), .O(n5356));
  invx  g04823(.a(n5356), .O(n5357));
  andx  g04824(.a(n4963), .b(n4956), .O(n5358));
  orx   g04825(.a(n5358), .b(n5357), .O(n5359));
  andx  g04826(.a(n5359), .b(n4961), .O(n5360));
  invx  g04827(.a(n5358), .O(n5361));
  andx  g04828(.a(n5361), .b(n5356), .O(n5362));
  andx  g04829(.a(n5362), .b(n4744), .O(n5363));
  orx   g04830(.a(n5363), .b(n5360), .O(n5364));
  andx  g04831(.a(n4490), .b(n403), .O(n5365));
  orx   g04832(.a(n5365), .b(n5354), .O(n5366));
  andx  g04833(.a(n5366), .b(n5364), .O(n5367));
  orx   g04834(.a(n5367), .b(n5355), .O(n5368));
  andx  g04835(.a(n4969), .b(n4974), .O(n5370));
  andx  g04836(.a(n4968), .b(n4966), .O(n5371));
  orx   g04837(.a(n5371), .b(n5370), .O(n5372));
  andx  g04838(.a(n5372), .b(n4738), .O(n5373));
  orx   g04839(.a(n4968), .b(n4966), .O(n5374));
  orx   g04840(.a(n4969), .b(n4974), .O(n5375));
  andx  g04841(.a(n5375), .b(n5374), .O(n5376));
  andx  g04842(.a(n5376), .b(n4971), .O(n5377));
  orx   g04843(.a(n5377), .b(n5373), .O(n5378));
  andx  g04844(.a(n5368), .b(n5378), .O(n5381));
  andx  g04845(.a(n5381), .b(n5088), .O(n5383));
  orx   g04846(.a(n5391), .b(n4720), .O(n5384));
  andx  g04847(.a(n5391), .b(n4720), .O(n5385));
  invx  g04848(.a(n5385), .O(n5386));
  andx  g04849(.a(n5386), .b(n5384), .O(n5387));
  invx  g04850(.a(n5387), .O(n5388));
  andx  g04851(.a(n5388), .b(n5383), .O(n5389));
  orx   g04852(.a(n5388), .b(n5383), .O(n5390));
  andx  g04853(.a(n5086), .b(n4728), .O(n5391));
  andx  g04854(.a(n5083), .b(n4727), .O(n5392));
  orx   g04855(.a(n5392), .b(n5391), .O(n5393));
  andx  g04856(.a(n5381), .b(n5393), .O(n5394));
  invx  g04857(.a(n5381), .O(n5395));
  andx  g04858(.a(n5395), .b(n5088), .O(n5396));
  orx   g04859(.a(n5396), .b(n5394), .O(n5397));
  invx  g04860(.a(n5368), .O(n5398));
  andx  g04861(.a(n5398), .b(n5378), .O(n5400));
  orx   g04862(.a(n5376), .b(n4971), .O(n5401));
  orx   g04863(.a(n5372), .b(n4738), .O(n5402));
  andx  g04864(.a(n5402), .b(n5401), .O(n5403));
  andx  g04865(.a(n5368), .b(n5403), .O(n5406));
  orx   g04866(.a(n5406), .b(n5400), .O(n5407));
  invx  g04867(.a(n5355), .O(n5408));
  andx  g04868(.a(n5366), .b(n5408), .O(n5409));
  orx   g04869(.a(n5409), .b(n5364), .O(n5410));
  orx   g04870(.a(n5362), .b(n4744), .O(n5411));
  orx   g04871(.a(n5359), .b(n4961), .O(n5412));
  andx  g04872(.a(n5412), .b(n5411), .O(n5413));
  invx  g04873(.a(n5409), .O(n5414));
  orx   g04874(.a(n5414), .b(n5413), .O(n5415));
  andx  g04875(.a(n5415), .b(n5410), .O(n5416));
  orx   g04876(.a(n5348), .b(n4950), .O(n5417));
  orx   g04877(.a(n5344), .b(n4752), .O(n5418));
  andx  g04878(.a(n5418), .b(n5417), .O(n5419));
  invx  g04879(.a(n5352), .O(n5420));
  orx   g04880(.a(n5420), .b(n5341), .O(n5421));
  andx  g04881(.a(n5421), .b(n5419), .O(n5422));
  invx  g04882(.a(n5341), .O(n5423));
  andx  g04883(.a(n5352), .b(n5423), .O(n5424));
  andx  g04884(.a(n5424), .b(n5350), .O(n5425));
  orx   g04885(.a(n5425), .b(n5422), .O(n5426));
  invx  g04886(.a(n5322), .O(n5427));
  invx  g04887(.a(n5323), .O(n5428));
  andx  g04888(.a(n5105), .b(n4925), .O(n5429));
  andx  g04889(.a(n5099), .b(n4915), .O(n5430));
  orx   g04890(.a(n5430), .b(n5429), .O(n5431));
  invx  g04891(.a(n5314), .O(n5432));
  andx  g04892(.a(n5432), .b(n5299), .O(n5433));
  andx  g04893(.a(n5432), .b(n5308), .O(n5434));
  orx   g04894(.a(n5434), .b(n5433), .O(n5435));
  orx   g04895(.a(n5435), .b(n5309), .O(n5436));
  andx  g04896(.a(n5436), .b(n5431), .O(n5437));
  orx   g04897(.a(n5437), .b(n5428), .O(n5438));
  andx  g04898(.a(n5438), .b(n5427), .O(n5439));
  orx   g04899(.a(n5439), .b(n4062), .O(n5440));
  andx  g04900(.a(n5338), .b(n5440), .O(n5441));
  orx   g04901(.a(n5441), .b(n5336), .O(n5442));
  orx   g04902(.a(n5334), .b(n4758), .O(n5443));
  orx   g04903(.a(n5330), .b(n4935), .O(n5444));
  andx  g04904(.a(n5444), .b(n5443), .O(n5445));
  invx  g04905(.a(n5337), .O(n5446));
  andx  g04906(.a(n5446), .b(n5439), .O(n5447));
  orx   g04907(.a(n5447), .b(n5327), .O(n5448));
  orx   g04908(.a(n5448), .b(n5445), .O(n5449));
  andx  g04909(.a(n5449), .b(n5442), .O(n5450));
  orx   g04910(.a(n5432), .b(n5299), .O(n5460));
  andx  g04911(.a(n5460), .b(n5315), .O(n5461));
  andx  g04912(.a(n5461), .b(n5318), .O(n5462));
  andx  g04913(.a(n5314), .b(n5313), .O(n5466));
  orx   g04914(.a(n5466), .b(n5433), .O(n5467));
  andx  g04915(.a(n5467), .b(n5308), .O(n5468));
  orx   g04916(.a(n5468), .b(n5462), .O(n5469));
  andx  g04917(.a(n5288), .b(n5296), .O(n5470));
  andx  g04918(.a(n5289), .b(n5286), .O(n5471));
  orx   g04919(.a(n5471), .b(n5470), .O(n5472));
  andx  g04920(.a(n5472), .b(n5139), .O(n5473));
  orx   g04921(.a(n5289), .b(n5286), .O(n5474));
  orx   g04922(.a(n5288), .b(n5296), .O(n5475));
  andx  g04923(.a(n5475), .b(n5474), .O(n5476));
  andx  g04924(.a(n5476), .b(n5293), .O(n5477));
  orx   g04925(.a(n5477), .b(n5473), .O(n5478));
  orx   g04926(.a(n5279), .b(n5249), .O(n5488));
  andx  g04927(.a(n5488), .b(n5265), .O(n5489));
  andx  g04928(.a(n5489), .b(n5268), .O(n5490));
  andx  g04929(.a(n5264), .b(n5263), .O(n5494));
  orx   g04930(.a(n5494), .b(n5280), .O(n5495));
  andx  g04931(.a(n5495), .b(n5258), .O(n5496));
  orx   g04932(.a(n5496), .b(n5490), .O(n5497));
  orx   g04933(.a(n5233), .b(n5231), .O(n5498));
  orx   g04934(.a(n5234), .b(n5217), .O(n5499));
  andx  g04935(.a(n5499), .b(n5498), .O(n5500));
  orx   g04936(.a(n5500), .b(n5170), .O(n5501));
  andx  g04937(.a(n5234), .b(n5217), .O(n5502));
  andx  g04938(.a(n5233), .b(n5231), .O(n5503));
  orx   g04939(.a(n5503), .b(n5502), .O(n5504));
  orx   g04940(.a(n5504), .b(n5222), .O(n5505));
  andx  g04941(.a(n5505), .b(n5501), .O(n5506));
  orx   g04942(.a(n5214), .b(n5228), .O(n5507));
  orx   g04943(.a(n5224), .b(n5212), .O(n5508));
  andx  g04944(.a(n5508), .b(n5507), .O(n5509));
  orx   g04945(.a(n5509), .b(n5227), .O(n5510));
  andx  g04946(.a(n5224), .b(n5212), .O(n5511));
  andx  g04947(.a(n5214), .b(n5228), .O(n5512));
  orx   g04948(.a(n5512), .b(n5511), .O(n5513));
  orx   g04949(.a(n5513), .b(n5179), .O(n5514));
  andx  g04950(.a(n5514), .b(n5510), .O(n5515));
  orx   g04951(.a(n3239), .b(n404), .O(n5516));
  orx   g04952(.a(n4790), .b(n5183), .O(n5517));
  orx   g04953(.a(n5181), .b(n4789), .O(n5518));
  andx  g04954(.a(n5518), .b(n5517), .O(n5519));
  orx   g04955(.a(n5519), .b(n5516), .O(n5520));
  invx  g04956(.a(n5189), .O(n5521));
  orx   g04957(.a(n5521), .b(n5516), .O(n5522));
  orx   g04958(.a(n5521), .b(n5519), .O(n5523));
  andx  g04959(.a(n5523), .b(n5522), .O(n5524));
  andx  g04960(.a(n5524), .b(n5520), .O(n5525));
  orx   g04961(.a(n3236), .b(n404), .O(n5526));
  andx  g04962(.a(n5526), .b(n5525), .O(n5527));
  orx   g04963(.a(n5527), .b(n5194), .O(n5528));
  andx  g04964(.a(n5528), .b(n5208), .O(n5529));
  andx  g04965(.a(n5201), .b(n5206), .O(n5530));
  andx  g04966(.a(n4787), .b(n5199), .O(n5531));
  orx   g04967(.a(n5531), .b(n5530), .O(n5532));
  orx   g04968(.a(n5525), .b(n3236), .O(n5533));
  andx  g04969(.a(n5210), .b(n5533), .O(n5534));
  andx  g04970(.a(n5534), .b(n5532), .O(n5535));
  orx   g04971(.a(n5535), .b(n5529), .O(n5536));
  andx  g04972(.a(n148), .b(pi04), .O(n5537));
  andx  g04973(.a(n153), .b(pi05), .O(n5538));
  andx  g04974(.a(n67), .b(pi02), .O(n5539));
  orx   g04975(.a(n5539), .b(n5538), .O(n5540));
  orx   g04976(.a(n5540), .b(n5537), .O(n5541));
  andx  g04977(.a(n159), .b(pi03), .O(n5542));
  andx  g04978(.a(n165), .b(pi06), .O(n5543));
  andx  g04979(.a(n161), .b(pi07), .O(n5544));
  andx  g04980(.a(n103), .b(pi08), .O(n5545));
  andx  g04981(.a(pi19), .b(pi09), .O(n5546));
  orx   g04982(.a(n5546), .b(n5545), .O(n5547));
  orx   g04983(.a(n5547), .b(n5544), .O(n5548));
  orx   g04984(.a(n5548), .b(n5543), .O(n5549));
  orx   g04985(.a(n5549), .b(n5542), .O(n5550));
  orx   g04986(.a(n5550), .b(n5541), .O(n5551));
  andx  g04987(.a(n5551), .b(n92), .O(n5552));
  andx  g04988(.a(n99), .b(pi01), .O(n5553));
  andx  g04989(.a(n143), .b(pi00), .O(n5554));
  orx   g04990(.a(n5554), .b(n5553), .O(n5555));
  orx   g04991(.a(n5555), .b(n5552), .O(n5556));
  andx  g04992(.a(n5556), .b(n3230), .O(n5557));
  invx  g04993(.a(n5188), .O(n5558));
  orx   g04994(.a(n5558), .b(n5187), .O(n5559));
  invx  g04995(.a(n5559), .O(n5560));
  andx  g04996(.a(n5558), .b(n5187), .O(n5561));
  orx   g04997(.a(n5561), .b(n5560), .O(n5562));
  andx  g04998(.a(n5562), .b(n5557), .O(n5563));
  andx  g04999(.a(n1790), .b(n403), .O(n5564));
  andx  g05000(.a(n5556), .b(n3258), .O(n5565));
  andx  g05001(.a(n5565), .b(n5564), .O(n5566));
  andx  g05002(.a(n5566), .b(n5557), .O(n5567));
  andx  g05003(.a(n5566), .b(n5562), .O(n5568));
  orx   g05004(.a(n5568), .b(n5567), .O(n5569));
  orx   g05005(.a(n5569), .b(n5563), .O(n5570));
  andx  g05006(.a(n5570), .b(n3221), .O(n5571));
  andx  g05007(.a(n5521), .b(n5180), .O(n5572));
  andx  g05008(.a(n5189), .b(n5516), .O(n5573));
  orx   g05009(.a(n5573), .b(n5572), .O(n5574));
  orx   g05010(.a(n5185), .b(n5574), .O(n5578));
  orx   g05011(.a(n5189), .b(n5516), .O(n5579));
  orx   g05012(.a(n5521), .b(n5180), .O(n5580));
  andx  g05013(.a(n5580), .b(n5579), .O(n5581));
  orx   g05014(.a(n5519), .b(n5581), .O(n5582));
  andx  g05015(.a(n5582), .b(n5578), .O(n5583));
  andx  g05016(.a(n5556), .b(n3221), .O(n5584));
  orx   g05017(.a(n5584), .b(n5570), .O(n5585));
  andx  g05018(.a(n5585), .b(n5583), .O(n5586));
  orx   g05019(.a(n5586), .b(n5571), .O(n5587));
  andx  g05020(.a(n5587), .b(n5536), .O(n5588));
  andx  g05021(.a(n5556), .b(n3210), .O(n5589));
  orx   g05022(.a(n5587), .b(n5536), .O(n5590));
  andx  g05023(.a(n5590), .b(n5589), .O(n5591));
  orx   g05024(.a(n5591), .b(n5588), .O(n5592));
  andx  g05025(.a(n5592), .b(n5515), .O(n5593));
  invx  g05026(.a(n5593), .O(n5594));
  andx  g05027(.a(n5513), .b(n5179), .O(n5595));
  andx  g05028(.a(n5509), .b(n5227), .O(n5596));
  orx   g05029(.a(n5596), .b(n5595), .O(n5597));
  orx   g05030(.a(n5534), .b(n5532), .O(n5598));
  orx   g05031(.a(n5528), .b(n5208), .O(n5599));
  andx  g05032(.a(n5599), .b(n5598), .O(n5600));
  invx  g05033(.a(n5563), .O(n5601));
  invx  g05034(.a(n5556), .O(n5602));
  orx   g05035(.a(n5602), .b(n3239), .O(n5603));
  invx  g05036(.a(n5566), .O(n5604));
  orx   g05037(.a(n5604), .b(n5603), .O(n5605));
  invx  g05038(.a(n5561), .O(n5606));
  andx  g05039(.a(n5606), .b(n5559), .O(n5607));
  orx   g05040(.a(n5604), .b(n5607), .O(n5608));
  andx  g05041(.a(n5608), .b(n5605), .O(n5609));
  andx  g05042(.a(n5609), .b(n5601), .O(n5610));
  orx   g05043(.a(n5610), .b(n3236), .O(n5611));
  andx  g05044(.a(n5519), .b(n5581), .O(n5612));
  andx  g05045(.a(n5185), .b(n5574), .O(n5613));
  orx   g05046(.a(n5613), .b(n5612), .O(n5614));
  orx   g05047(.a(n5602), .b(n3236), .O(n5615));
  andx  g05048(.a(n5615), .b(n5610), .O(n5616));
  orx   g05049(.a(n5616), .b(n5614), .O(n5617));
  andx  g05050(.a(n5617), .b(n5611), .O(n5618));
  orx   g05051(.a(n5618), .b(n5600), .O(n5619));
  orx   g05052(.a(n5602), .b(n3270), .O(n5620));
  andx  g05053(.a(n5618), .b(n5600), .O(n5621));
  orx   g05054(.a(n5621), .b(n5620), .O(n5622));
  andx  g05055(.a(n5622), .b(n5619), .O(n5623));
  andx  g05056(.a(n5623), .b(n5597), .O(n5624));
  orx   g05057(.a(n5602), .b(n3201), .O(n5625));
  orx   g05058(.a(n5625), .b(n5624), .O(n5626));
  andx  g05059(.a(n5626), .b(n5594), .O(n5627));
  andx  g05060(.a(n5627), .b(n5506), .O(n5628));
  andx  g05061(.a(n5556), .b(n3180), .O(n5629));
  invx  g05062(.a(n5629), .O(n5630));
  orx   g05063(.a(n5630), .b(n5628), .O(n5631));
  andx  g05064(.a(n5504), .b(n5222), .O(n5632));
  andx  g05065(.a(n5500), .b(n5170), .O(n5633));
  orx   g05066(.a(n5633), .b(n5632), .O(n5634));
  orx   g05067(.a(n5592), .b(n5515), .O(n5635));
  andx  g05068(.a(n5556), .b(n3284), .O(n5636));
  andx  g05069(.a(n5636), .b(n5635), .O(n5637));
  orx   g05070(.a(n5637), .b(n5593), .O(n5638));
  andx  g05071(.a(n5638), .b(n5634), .O(n5639));
  invx  g05072(.a(n5639), .O(n5640));
  andx  g05073(.a(n5640), .b(n5631), .O(n5641));
  andx  g05074(.a(n5239), .b(n5236), .O(n5642));
  andx  g05075(.a(n5238), .b(n5246), .O(n5643));
  orx   g05076(.a(n5643), .b(n5642), .O(n5644));
  andx  g05077(.a(n5644), .b(n5161), .O(n5645));
  orx   g05078(.a(n5238), .b(n5246), .O(n5646));
  orx   g05079(.a(n5239), .b(n5236), .O(n5647));
  andx  g05080(.a(n5647), .b(n5646), .O(n5648));
  andx  g05081(.a(n5648), .b(n5243), .O(n5649));
  orx   g05082(.a(n5649), .b(n5645), .O(n5650));
  andx  g05083(.a(n5650), .b(n5641), .O(n5651));
  andx  g05084(.a(n5556), .b(n3429), .O(n5652));
  invx  g05085(.a(n5652), .O(n5653));
  andx  g05086(.a(n5653), .b(n5641), .O(n5654));
  andx  g05087(.a(n5653), .b(n5650), .O(n5655));
  orx   g05088(.a(n5655), .b(n5654), .O(n5656));
  orx   g05089(.a(n5656), .b(n5651), .O(n5657));
  andx  g05090(.a(n5657), .b(n5497), .O(n5658));
  andx  g05091(.a(n5556), .b(n3171), .O(n5659));
  invx  g05092(.a(n5659), .O(n5660));
  orx   g05093(.a(n5660), .b(n5658), .O(n5661));
  orx   g05094(.a(n5495), .b(n5258), .O(n5662));
  orx   g05095(.a(n5489), .b(n5268), .O(n5663));
  andx  g05096(.a(n5663), .b(n5662), .O(n5664));
  invx  g05097(.a(n5651), .O(n5665));
  orx   g05098(.a(n5638), .b(n5634), .O(n5666));
  andx  g05099(.a(n5629), .b(n5666), .O(n5667));
  orx   g05100(.a(n5639), .b(n5667), .O(n5668));
  orx   g05101(.a(n5652), .b(n5668), .O(n5669));
  orx   g05102(.a(n5648), .b(n5243), .O(n5670));
  orx   g05103(.a(n5644), .b(n5161), .O(n5671));
  andx  g05104(.a(n5671), .b(n5670), .O(n5672));
  orx   g05105(.a(n5652), .b(n5672), .O(n5673));
  andx  g05106(.a(n5673), .b(n5669), .O(n5674));
  andx  g05107(.a(n5674), .b(n5665), .O(n5675));
  andx  g05108(.a(n5675), .b(n5664), .O(n5676));
  invx  g05109(.a(n5676), .O(n5677));
  andx  g05110(.a(n5677), .b(n5661), .O(n5678));
  andx  g05111(.a(n5275), .b(n5283), .O(n5679));
  andx  g05112(.a(n5274), .b(n5271), .O(n5680));
  orx   g05113(.a(n5680), .b(n5679), .O(n5681));
  andx  g05114(.a(n5681), .b(n5278), .O(n5682));
  orx   g05115(.a(n5274), .b(n5271), .O(n5683));
  orx   g05116(.a(n5275), .b(n5283), .O(n5684));
  andx  g05117(.a(n5684), .b(n5683), .O(n5685));
  andx  g05118(.a(n5685), .b(n5152), .O(n5686));
  orx   g05119(.a(n5686), .b(n5682), .O(n5687));
  andx  g05120(.a(n5687), .b(n5678), .O(n5688));
  andx  g05121(.a(n5556), .b(n3413), .O(n5689));
  invx  g05122(.a(n5689), .O(n5690));
  andx  g05123(.a(n5690), .b(n5678), .O(n5691));
  andx  g05124(.a(n5690), .b(n5687), .O(n5692));
  orx   g05125(.a(n5692), .b(n5691), .O(n5693));
  orx   g05126(.a(n5693), .b(n5688), .O(n5694));
  andx  g05127(.a(n5694), .b(n5478), .O(n5695));
  andx  g05128(.a(n5556), .b(n3645), .O(n5696));
  invx  g05129(.a(n5696), .O(n5697));
  andx  g05130(.a(n5697), .b(n5478), .O(n5698));
  andx  g05131(.a(n5697), .b(n5694), .O(n5699));
  orx   g05132(.a(n5699), .b(n5698), .O(n5700));
  orx   g05133(.a(n5700), .b(n5695), .O(n5701));
  andx  g05134(.a(n5701), .b(n5469), .O(n5702));
  andx  g05135(.a(n5556), .b(n3721), .O(n5703));
  invx  g05136(.a(n5703), .O(n5704));
  orx   g05137(.a(n5704), .b(n5702), .O(n5705));
  orx   g05138(.a(n5467), .b(n5308), .O(n5706));
  orx   g05139(.a(n5461), .b(n5318), .O(n5707));
  andx  g05140(.a(n5707), .b(n5706), .O(n5708));
  invx  g05141(.a(n5695), .O(n5709));
  orx   g05142(.a(n5476), .b(n5293), .O(n5710));
  orx   g05143(.a(n5472), .b(n5139), .O(n5711));
  andx  g05144(.a(n5711), .b(n5710), .O(n5712));
  orx   g05145(.a(n5696), .b(n5712), .O(n5713));
  invx  g05146(.a(n5699), .O(n5714));
  andx  g05147(.a(n5714), .b(n5713), .O(n5715));
  andx  g05148(.a(n5715), .b(n5709), .O(n5716));
  andx  g05149(.a(n5716), .b(n5708), .O(n5717));
  invx  g05150(.a(n5717), .O(n5718));
  andx  g05151(.a(n5718), .b(n5705), .O(n5719));
  orx   g05152(.a(n5323), .b(n5436), .O(n5720));
  orx   g05153(.a(n5428), .b(n5321), .O(n5721));
  andx  g05154(.a(n5721), .b(n5720), .O(n5722));
  andx  g05155(.a(n5722), .b(n5431), .O(n5723));
  andx  g05156(.a(n5428), .b(n5321), .O(n5724));
  andx  g05157(.a(n5323), .b(n5436), .O(n5725));
  orx   g05158(.a(n5725), .b(n5724), .O(n5726));
  andx  g05159(.a(n5726), .b(n5107), .O(n5727));
  orx   g05160(.a(n5727), .b(n5723), .O(n5728));
  andx  g05161(.a(n5728), .b(n5719), .O(n5729));
  invx  g05162(.a(n5729), .O(n5730));
  orx   g05163(.a(n5716), .b(n5708), .O(n5731));
  andx  g05164(.a(n5703), .b(n5731), .O(n5732));
  orx   g05165(.a(n5717), .b(n5732), .O(n5733));
  andx  g05166(.a(n5556), .b(n4063), .O(n5734));
  orx   g05167(.a(n5734), .b(n5733), .O(n5735));
  orx   g05168(.a(n5726), .b(n5107), .O(n5736));
  orx   g05169(.a(n5722), .b(n5431), .O(n5737));
  andx  g05170(.a(n5737), .b(n5736), .O(n5738));
  orx   g05171(.a(n5734), .b(n5738), .O(n5739));
  andx  g05172(.a(n5739), .b(n5735), .O(n5740));
  andx  g05173(.a(n5740), .b(n5730), .O(n5741));
  andx  g05174(.a(n5741), .b(n5450), .O(n5742));
  invx  g05175(.a(n5742), .O(n5743));
  andx  g05176(.a(n5448), .b(n5445), .O(n5744));
  andx  g05177(.a(n5441), .b(n5336), .O(n5745));
  orx   g05178(.a(n5745), .b(n5744), .O(n5746));
  invx  g05179(.a(n5734), .O(n5747));
  andx  g05180(.a(n5747), .b(n5719), .O(n5748));
  andx  g05181(.a(n5747), .b(n5728), .O(n5749));
  orx   g05182(.a(n5749), .b(n5748), .O(n5750));
  orx   g05183(.a(n5750), .b(n5729), .O(n5751));
  andx  g05184(.a(n5751), .b(n5746), .O(n5752));
  andx  g05185(.a(n5556), .b(n4114), .O(n5753));
  invx  g05186(.a(n5753), .O(n5754));
  orx   g05187(.a(n5754), .b(n5752), .O(n5755));
  andx  g05188(.a(n5755), .b(n5743), .O(n5756));
  andx  g05189(.a(n5756), .b(n5426), .O(n5757));
  andx  g05190(.a(n5556), .b(n4490), .O(n5758));
  invx  g05191(.a(n5758), .O(n5759));
  orx   g05192(.a(n5759), .b(n5757), .O(n5760));
  orx   g05193(.a(n5424), .b(n5350), .O(n5761));
  orx   g05194(.a(n5421), .b(n5419), .O(n5762));
  andx  g05195(.a(n5762), .b(n5761), .O(n5763));
  orx   g05196(.a(n5741), .b(n5450), .O(n5764));
  andx  g05197(.a(n5753), .b(n5764), .O(n5765));
  orx   g05198(.a(n5765), .b(n5742), .O(n5766));
  andx  g05199(.a(n5766), .b(n5763), .O(n5767));
  invx  g05200(.a(n5767), .O(n5768));
  andx  g05201(.a(n5768), .b(n5760), .O(n5769));
  invx  g05202(.a(n5769), .O(n5770));
  andx  g05203(.a(n5770), .b(n5416), .O(n5771));
  andx  g05204(.a(n5556), .b(n2724), .O(n5772));
  andx  g05205(.a(n5771), .b(n5407), .O(n5777));
  andx  g05206(.a(n5777), .b(n5397), .O(n5778));
  andx  g05207(.a(n5778), .b(n5390), .O(n5779));
  orx   g05208(.a(n5779), .b(n5389), .O(n5780));
  orx   g05209(.a(n5076), .b(n4983), .O(n5781));
  andx  g05210(.a(n5781), .b(n5780), .O(n5782));
  orx   g05211(.a(n5782), .b(n5079), .O(n5783));
  invx  g05212(.a(n5005), .O(n5784));
  andx  g05213(.a(n5011), .b(n5784), .O(n5785));
  invx  g05214(.a(n5785), .O(n5786));
  andx  g05215(.a(n5010), .b(n5005), .O(n5787));
  orx   g05216(.a(n5787), .b(n5013), .O(n5788));
  andx  g05217(.a(n5788), .b(n5786), .O(n5789));
  andx  g05218(.a(n4063), .b(n299), .O(n5790));
  andx  g05219(.a(n5790), .b(n5789), .O(n5791));
  invx  g05220(.a(n5789), .O(n5792));
  invx  g05221(.a(n5790), .O(n5793));
  andx  g05222(.a(n5793), .b(n5792), .O(n5794));
  orx   g05223(.a(n5794), .b(n5791), .O(n5795));
  andx  g05224(.a(n4509), .b(n827), .O(n5796));
  andx  g05225(.a(n5796), .b(n3721), .O(n5797));
  andx  g05226(.a(n3721), .b(n827), .O(n5798));
  invx  g05227(.a(n5798), .O(n5799));
  andx  g05228(.a(n5799), .b(n3645), .O(n5800));
  orx   g05229(.a(n5800), .b(n5797), .O(n5801));
  andx  g05230(.a(n5001), .b(n3415), .O(n5802));
  orx   g05231(.a(n5802), .b(n4509), .O(n5803));
  andx  g05232(.a(n5000), .b(n5803), .O(n5806));
  andx  g05233(.a(n5806), .b(n5801), .O(n5807));
  invx  g05234(.a(n5807), .O(n5808));
  orx   g05235(.a(n5806), .b(n5801), .O(n5809));
  andx  g05236(.a(n5809), .b(n5808), .O(n5810));
  invx  g05237(.a(n5810), .O(n5811));
  andx  g05238(.a(n5811), .b(n5795), .O(n5812));
  invx  g05239(.a(n5812), .O(n5813));
  orx   g05240(.a(n5811), .b(n5795), .O(n5814));
  andx  g05241(.a(n5814), .b(n5813), .O(n5815));
  invx  g05242(.a(n5815), .O(n5816));
  andx  g05243(.a(n5026), .b(n5030), .O(n5817));
  orx   g05244(.a(n5817), .b(n5023), .O(n5818));
  andx  g05245(.a(n5818), .b(n4114), .O(n5819));
  invx  g05246(.a(n5819), .O(n5820));
  andx  g05247(.a(n4114), .b(n338), .O(n5821));
  orx   g05248(.a(n5821), .b(n5818), .O(n5822));
  andx  g05249(.a(n5822), .b(n5820), .O(n5823));
  invx  g05250(.a(n5823), .O(n5824));
  andx  g05251(.a(n5824), .b(n5816), .O(n5825));
  andx  g05252(.a(n5823), .b(n5815), .O(n5826));
  orx   g05253(.a(n5826), .b(n5825), .O(n5827));
  invx  g05254(.a(n5032), .O(n5830));
  andx  g05255(.a(n5037), .b(n5830), .O(n5831));
  invx  g05256(.a(n5831), .O(n5832));
  andx  g05257(.a(n5036), .b(n5032), .O(n5833));
  orx   g05258(.a(n5833), .b(n5039), .O(n5834));
  andx  g05259(.a(n5834), .b(n5832), .O(n5835));
  andx  g05260(.a(n5835), .b(n376), .O(n5838));
  andx  g05261(.a(n5838), .b(n5827), .O(n5840));
  invx  g05262(.a(n5840), .O(n5841));
  orx   g05263(.a(n5838), .b(n5827), .O(n5842));
  andx  g05264(.a(n5842), .b(n5841), .O(n5843));
  andx  g05265(.a(n5052), .b(n5056), .O(n5844));
  orx   g05266(.a(n5844), .b(n5049), .O(n5845));
  andx  g05267(.a(n5845), .b(n2724), .O(n5846));
  invx  g05268(.a(n5845), .O(n5851));
  andx  g05269(.a(n5851), .b(n5843), .O(n5852));
  invx  g05270(.a(n5843), .O(n5853));
  orx   g05271(.a(n7660), .b(n5852), .O(n5855));
  invx  g05272(.a(n5058), .O(n5856));
  andx  g05273(.a(n5065), .b(n5856), .O(n5858));
  andx  g05274(.a(n5858), .b(n5855), .O(n5862));
  invx  g05275(.a(n5855), .O(n5863));
  invx  g05276(.a(n5858), .O(n5864));
  andx  g05277(.a(n5864), .b(n5863), .O(n5865));
  orx   g05278(.a(n5865), .b(n5862), .O(n5866));
  andx  g05279(.a(n5866), .b(n5783), .O(n5867));
  andx  g05280(.a(n5759), .b(n5766), .O(n5868));
  andx  g05281(.a(n5758), .b(n5756), .O(n5869));
  orx   g05282(.a(n5869), .b(n5868), .O(n5870));
  andx  g05283(.a(n5870), .b(n5426), .O(n5871));
  orx   g05284(.a(n5758), .b(n5756), .O(n5872));
  orx   g05285(.a(n5759), .b(n5766), .O(n5873));
  andx  g05286(.a(n5873), .b(n5872), .O(n5874));
  andx  g05287(.a(n5874), .b(n5763), .O(n5875));
  orx   g05288(.a(n5875), .b(n5871), .O(n5876));
  invx  g05289(.a(n4490), .O(n5878));
  andx  g05290(.a(n5734), .b(n5733), .O(n5888));
  orx   g05291(.a(n5888), .b(n5748), .O(n5889));
  orx   g05292(.a(n5889), .b(n5728), .O(n5890));
  orx   g05293(.a(n5747), .b(n5719), .O(n5894));
  andx  g05294(.a(n5894), .b(n5735), .O(n5895));
  orx   g05295(.a(n5895), .b(n5738), .O(n5896));
  andx  g05296(.a(n5896), .b(n5890), .O(n5897));
  orx   g05297(.a(n5689), .b(n5678), .O(n5901));
  orx   g05298(.a(n5675), .b(n5664), .O(n5902));
  andx  g05299(.a(n5659), .b(n5902), .O(n5903));
  orx   g05300(.a(n5676), .b(n5903), .O(n5904));
  orx   g05301(.a(n5690), .b(n5904), .O(n5905));
  andx  g05302(.a(n5905), .b(n5901), .O(n5906));
  orx   g05303(.a(n5906), .b(n5687), .O(n5907));
  andx  g05304(.a(n5685), .b(n5278), .O(n5908));
  andx  g05305(.a(n5681), .b(n5152), .O(n5909));
  orx   g05306(.a(n5909), .b(n5908), .O(n5910));
  andx  g05307(.a(n5690), .b(n5904), .O(n5911));
  andx  g05308(.a(n5689), .b(n5678), .O(n5912));
  orx   g05309(.a(n5912), .b(n5911), .O(n5913));
  orx   g05310(.a(n5913), .b(n5910), .O(n5914));
  andx  g05311(.a(n5914), .b(n5907), .O(n5915));
  orx   g05312(.a(n5589), .b(n5618), .O(n5916));
  orx   g05313(.a(n5620), .b(n5587), .O(n5917));
  andx  g05314(.a(n5917), .b(n5916), .O(n5918));
  orx   g05315(.a(n5918), .b(n5600), .O(n5919));
  andx  g05316(.a(n5620), .b(n5587), .O(n5920));
  andx  g05317(.a(n5589), .b(n5618), .O(n5921));
  orx   g05318(.a(n5921), .b(n5920), .O(n5922));
  orx   g05319(.a(n5922), .b(n5536), .O(n5923));
  andx  g05320(.a(n5923), .b(n5919), .O(n5924));
  orx   g05321(.a(n5616), .b(n5571), .O(n5925));
  andx  g05322(.a(n5925), .b(n5583), .O(n5926));
  andx  g05323(.a(n5585), .b(n5611), .O(n5927));
  andx  g05324(.a(n5927), .b(n5614), .O(n5928));
  orx   g05325(.a(n5928), .b(n5926), .O(n5929));
  andx  g05326(.a(n99), .b(pi00), .O(n5930));
  andx  g05327(.a(n148), .b(pi03), .O(n5931));
  andx  g05328(.a(n67), .b(pi01), .O(n5932));
  andx  g05329(.a(n153), .b(pi04), .O(n5933));
  orx   g05330(.a(n5933), .b(n5932), .O(n5934));
  orx   g05331(.a(n5934), .b(n5931), .O(n5935));
  andx  g05332(.a(n159), .b(pi02), .O(n5936));
  andx  g05333(.a(n161), .b(pi06), .O(n5937));
  andx  g05334(.a(n165), .b(pi05), .O(n5938));
  andx  g05335(.a(pi19), .b(pi08), .O(n5939));
  andx  g05336(.a(n103), .b(pi07), .O(n5940));
  orx   g05337(.a(n5940), .b(n5939), .O(n5941));
  orx   g05338(.a(n5941), .b(n5938), .O(n5942));
  orx   g05339(.a(n5942), .b(n5937), .O(n5943));
  orx   g05340(.a(n5943), .b(n5936), .O(n5944));
  orx   g05341(.a(n5944), .b(n5935), .O(n5945));
  andx  g05342(.a(n5945), .b(n92), .O(n5946));
  orx   g05343(.a(n5946), .b(n5930), .O(n5947));
  andx  g05344(.a(n5947), .b(n3230), .O(n5948));
  invx  g05345(.a(n5565), .O(n5949));
  andx  g05346(.a(n5949), .b(n5564), .O(n5950));
  invx  g05347(.a(n5564), .O(n5951));
  andx  g05348(.a(n5565), .b(n5951), .O(n5952));
  orx   g05349(.a(n5952), .b(n5950), .O(n5953));
  andx  g05350(.a(n5953), .b(n5948), .O(n5954));
  andx  g05351(.a(n5556), .b(n1790), .O(n5955));
  andx  g05352(.a(n5947), .b(n3258), .O(n5956));
  andx  g05353(.a(n5956), .b(n5955), .O(n5957));
  andx  g05354(.a(n5957), .b(n5948), .O(n5958));
  andx  g05355(.a(n5957), .b(n5953), .O(n5959));
  orx   g05356(.a(n5959), .b(n5958), .O(n5960));
  orx   g05357(.a(n5960), .b(n5954), .O(n5961));
  andx  g05358(.a(n5961), .b(n3221), .O(n5962));
  andx  g05359(.a(n5604), .b(n5557), .O(n5963));
  andx  g05360(.a(n5566), .b(n5603), .O(n5964));
  orx   g05361(.a(n5964), .b(n5963), .O(n5965));
  orx   g05362(.a(n5562), .b(n5965), .O(n5970));
  andx  g05363(.a(n5562), .b(n5965), .O(n5971));
  invx  g05364(.a(n5971), .O(n5972));
  andx  g05365(.a(n5972), .b(n5970), .O(n5973));
  andx  g05366(.a(n5947), .b(n3221), .O(n5974));
  orx   g05367(.a(n5974), .b(n5961), .O(n5975));
  andx  g05368(.a(n5975), .b(n5973), .O(n5976));
  orx   g05369(.a(n5976), .b(n5962), .O(n5977));
  andx  g05370(.a(n5977), .b(n5929), .O(n5978));
  andx  g05371(.a(n5947), .b(n3210), .O(n5979));
  orx   g05372(.a(n5977), .b(n5929), .O(n5980));
  andx  g05373(.a(n5980), .b(n5979), .O(n5981));
  orx   g05374(.a(n5981), .b(n5978), .O(n5982));
  andx  g05375(.a(n5982), .b(n5924), .O(n5983));
  invx  g05376(.a(n5983), .O(n5984));
  andx  g05377(.a(n5922), .b(n5536), .O(n5985));
  andx  g05378(.a(n5918), .b(n5600), .O(n5986));
  orx   g05379(.a(n5986), .b(n5985), .O(n5987));
  invx  g05380(.a(n5978), .O(n5988));
  invx  g05381(.a(n5979), .O(n5989));
  orx   g05382(.a(n5927), .b(n5614), .O(n5990));
  orx   g05383(.a(n5925), .b(n5583), .O(n5991));
  andx  g05384(.a(n5991), .b(n5990), .O(n5992));
  invx  g05385(.a(n5962), .O(n5993));
  invx  g05386(.a(n5970), .O(n5994));
  orx   g05387(.a(n5971), .b(n5994), .O(n5995));
  invx  g05388(.a(n5975), .O(n5996));
  orx   g05389(.a(n5996), .b(n5995), .O(n5997));
  andx  g05390(.a(n5997), .b(n5993), .O(n5998));
  andx  g05391(.a(n5998), .b(n5992), .O(n5999));
  orx   g05392(.a(n5999), .b(n5989), .O(n6000));
  andx  g05393(.a(n6000), .b(n5988), .O(n6001));
  andx  g05394(.a(n6001), .b(n5987), .O(n6002));
  invx  g05395(.a(n5947), .O(n6003));
  orx   g05396(.a(n6003), .b(n3201), .O(n6004));
  orx   g05397(.a(n6004), .b(n6002), .O(n6005));
  andx  g05398(.a(n6005), .b(n5984), .O(n6006));
  orx   g05399(.a(n5636), .b(n5623), .O(n6007));
  orx   g05400(.a(n5625), .b(n5592), .O(n6008));
  andx  g05401(.a(n6008), .b(n6007), .O(n6009));
  orx   g05402(.a(n6009), .b(n5515), .O(n6010));
  andx  g05403(.a(n5625), .b(n5592), .O(n6011));
  andx  g05404(.a(n5636), .b(n5623), .O(n6012));
  orx   g05405(.a(n6012), .b(n6011), .O(n6013));
  orx   g05406(.a(n6013), .b(n5597), .O(n6014));
  andx  g05407(.a(n6014), .b(n6010), .O(n6015));
  andx  g05408(.a(n6015), .b(n6006), .O(n6016));
  orx   g05409(.a(n6003), .b(n3183), .O(n6017));
  orx   g05410(.a(n6017), .b(n6016), .O(n6018));
  orx   g05411(.a(n6015), .b(n6006), .O(n6019));
  andx  g05412(.a(n6019), .b(n6018), .O(n6020));
  andx  g05413(.a(n5630), .b(n5627), .O(n6021));
  andx  g05414(.a(n5629), .b(n5638), .O(n6022));
  orx   g05415(.a(n6022), .b(n6021), .O(n6023));
  andx  g05416(.a(n6023), .b(n5506), .O(n6024));
  orx   g05417(.a(n5629), .b(n5638), .O(n6025));
  orx   g05418(.a(n5630), .b(n5627), .O(n6026));
  andx  g05419(.a(n6026), .b(n6025), .O(n6027));
  andx  g05420(.a(n6027), .b(n5634), .O(n6028));
  orx   g05421(.a(n6028), .b(n6024), .O(n6029));
  andx  g05422(.a(n6029), .b(n6020), .O(n6030));
  orx   g05423(.a(n6003), .b(n3297), .O(n6031));
  andx  g05424(.a(n6031), .b(n6020), .O(n6032));
  andx  g05425(.a(n6031), .b(n6029), .O(n6033));
  orx   g05426(.a(n6033), .b(n6032), .O(n6034));
  orx   g05427(.a(n6034), .b(n6030), .O(n6035));
  orx   g05428(.a(n5653), .b(n5641), .O(n6045));
  andx  g05429(.a(n6045), .b(n5669), .O(n6046));
  andx  g05430(.a(n6046), .b(n5672), .O(n6047));
  andx  g05431(.a(n5652), .b(n5668), .O(n6051));
  orx   g05432(.a(n6051), .b(n5654), .O(n6052));
  andx  g05433(.a(n6052), .b(n5650), .O(n6053));
  orx   g05434(.a(n6053), .b(n6047), .O(n6054));
  andx  g05435(.a(n6054), .b(n6035), .O(n6055));
  andx  g05436(.a(n5947), .b(n3171), .O(n6056));
  invx  g05437(.a(n6056), .O(n6057));
  orx   g05438(.a(n6057), .b(n6055), .O(n6058));
  invx  g05439(.a(n6030), .O(n6059));
  orx   g05440(.a(n5982), .b(n5924), .O(n6060));
  andx  g05441(.a(n5947), .b(n3284), .O(n6061));
  andx  g05442(.a(n6061), .b(n6060), .O(n6062));
  orx   g05443(.a(n6062), .b(n5983), .O(n6063));
  andx  g05444(.a(n6013), .b(n5597), .O(n6064));
  andx  g05445(.a(n6009), .b(n5515), .O(n6065));
  orx   g05446(.a(n6065), .b(n6064), .O(n6066));
  orx   g05447(.a(n6066), .b(n6063), .O(n6067));
  andx  g05448(.a(n5947), .b(n3180), .O(n6068));
  andx  g05449(.a(n6068), .b(n6067), .O(n6069));
  andx  g05450(.a(n6066), .b(n6063), .O(n6070));
  orx   g05451(.a(n6070), .b(n6069), .O(n6071));
  andx  g05452(.a(n5947), .b(n3429), .O(n6072));
  orx   g05453(.a(n6072), .b(n6071), .O(n6073));
  orx   g05454(.a(n6027), .b(n5634), .O(n6074));
  orx   g05455(.a(n6023), .b(n5506), .O(n6075));
  andx  g05456(.a(n6075), .b(n6074), .O(n6076));
  orx   g05457(.a(n6072), .b(n6076), .O(n6077));
  andx  g05458(.a(n6077), .b(n6073), .O(n6078));
  andx  g05459(.a(n6078), .b(n6059), .O(n6079));
  orx   g05460(.a(n6052), .b(n5650), .O(n6080));
  orx   g05461(.a(n6046), .b(n5672), .O(n6081));
  andx  g05462(.a(n6081), .b(n6080), .O(n6082));
  andx  g05463(.a(n6082), .b(n6079), .O(n6083));
  invx  g05464(.a(n6083), .O(n6084));
  andx  g05465(.a(n6084), .b(n6058), .O(n6085));
  orx   g05466(.a(n5659), .b(n5657), .O(n6086));
  orx   g05467(.a(n5660), .b(n5675), .O(n6087));
  andx  g05468(.a(n6087), .b(n6086), .O(n6088));
  andx  g05469(.a(n6088), .b(n5497), .O(n6089));
  andx  g05470(.a(n5660), .b(n5675), .O(n6090));
  andx  g05471(.a(n5659), .b(n5657), .O(n6091));
  orx   g05472(.a(n6091), .b(n6090), .O(n6092));
  andx  g05473(.a(n6092), .b(n5664), .O(n6093));
  orx   g05474(.a(n6093), .b(n6089), .O(n6094));
  andx  g05475(.a(n6094), .b(n6085), .O(n6095));
  invx  g05476(.a(n6095), .O(n6096));
  orx   g05477(.a(n6082), .b(n6079), .O(n6097));
  andx  g05478(.a(n6056), .b(n6097), .O(n6098));
  orx   g05479(.a(n6083), .b(n6098), .O(n6099));
  andx  g05480(.a(n5947), .b(n3413), .O(n6100));
  orx   g05481(.a(n6100), .b(n6099), .O(n6101));
  orx   g05482(.a(n6092), .b(n5664), .O(n6102));
  orx   g05483(.a(n6088), .b(n5497), .O(n6103));
  andx  g05484(.a(n6103), .b(n6102), .O(n6104));
  orx   g05485(.a(n6100), .b(n6104), .O(n6105));
  andx  g05486(.a(n6105), .b(n6101), .O(n6106));
  andx  g05487(.a(n6106), .b(n6096), .O(n6107));
  andx  g05488(.a(n6107), .b(n5915), .O(n6108));
  invx  g05489(.a(n6108), .O(n6109));
  andx  g05490(.a(n5947), .b(n3645), .O(n6110));
  invx  g05491(.a(n6110), .O(n6111));
  andx  g05492(.a(n5913), .b(n5910), .O(n6112));
  andx  g05493(.a(n5906), .b(n5687), .O(n6113));
  orx   g05494(.a(n6113), .b(n6112), .O(n6114));
  invx  g05495(.a(n6100), .O(n6115));
  andx  g05496(.a(n6115), .b(n6085), .O(n6116));
  andx  g05497(.a(n6115), .b(n6094), .O(n6117));
  orx   g05498(.a(n6117), .b(n6116), .O(n6118));
  orx   g05499(.a(n6118), .b(n6095), .O(n6119));
  andx  g05500(.a(n6119), .b(n6114), .O(n6120));
  orx   g05501(.a(n6120), .b(n6111), .O(n6121));
  andx  g05502(.a(n6121), .b(n6109), .O(n6122));
  andx  g05503(.a(n5696), .b(n5694), .O(n6123));
  invx  g05504(.a(n5688), .O(n6124));
  invx  g05505(.a(n5691), .O(n6125));
  orx   g05506(.a(n5689), .b(n5910), .O(n6129));
  andx  g05507(.a(n6129), .b(n6125), .O(n6130));
  andx  g05508(.a(n6130), .b(n6124), .O(n6131));
  andx  g05509(.a(n5697), .b(n6131), .O(n6132));
  orx   g05510(.a(n6132), .b(n6123), .O(n6133));
  andx  g05511(.a(n5712), .b(n6133), .O(n6143));
  orx   g05512(.a(n5697), .b(n6131), .O(n6144));
  orx   g05513(.a(n5696), .b(n5694), .O(n6145));
  andx  g05514(.a(n6145), .b(n6144), .O(n6146));
  andx  g05515(.a(n5478), .b(n6146), .O(n6150));
  orx   g05516(.a(n6150), .b(n6143), .O(n6151));
  andx  g05517(.a(n6151), .b(n6122), .O(n6152));
  andx  g05518(.a(n5947), .b(n3721), .O(n6153));
  invx  g05519(.a(n6153), .O(n6154));
  orx   g05520(.a(n6154), .b(n6152), .O(n6155));
  orx   g05521(.a(n6107), .b(n5915), .O(n6156));
  andx  g05522(.a(n6156), .b(n6110), .O(n6157));
  orx   g05523(.a(n6157), .b(n6108), .O(n6158));
  orx   g05524(.a(n5478), .b(n6146), .O(n6159));
  orx   g05525(.a(n5712), .b(n6133), .O(n6160));
  andx  g05526(.a(n6160), .b(n6159), .O(n6161));
  andx  g05527(.a(n6161), .b(n6158), .O(n6162));
  invx  g05528(.a(n6162), .O(n6163));
  andx  g05529(.a(n6163), .b(n6155), .O(n6164));
  orx   g05530(.a(n5703), .b(n5701), .O(n6165));
  orx   g05531(.a(n5704), .b(n5716), .O(n6166));
  andx  g05532(.a(n6166), .b(n6165), .O(n6167));
  andx  g05533(.a(n6167), .b(n5469), .O(n6168));
  andx  g05534(.a(n5704), .b(n5716), .O(n6169));
  andx  g05535(.a(n5703), .b(n5701), .O(n6170));
  orx   g05536(.a(n6170), .b(n6169), .O(n6171));
  andx  g05537(.a(n6171), .b(n5708), .O(n6172));
  orx   g05538(.a(n6172), .b(n6168), .O(n6173));
  andx  g05539(.a(n6173), .b(n6164), .O(n6174));
  invx  g05540(.a(n6174), .O(n6175));
  orx   g05541(.a(n6161), .b(n6158), .O(n6176));
  andx  g05542(.a(n6153), .b(n6176), .O(n6177));
  orx   g05543(.a(n6162), .b(n6177), .O(n6178));
  andx  g05544(.a(n5947), .b(n4063), .O(n6179));
  orx   g05545(.a(n6179), .b(n6178), .O(n6180));
  orx   g05546(.a(n6171), .b(n5708), .O(n6181));
  orx   g05547(.a(n6167), .b(n5469), .O(n6182));
  andx  g05548(.a(n6182), .b(n6181), .O(n6183));
  orx   g05549(.a(n6179), .b(n6183), .O(n6184));
  andx  g05550(.a(n6184), .b(n6180), .O(n6185));
  andx  g05551(.a(n6185), .b(n6175), .O(n6186));
  andx  g05552(.a(n6186), .b(n5897), .O(n6187));
  invx  g05553(.a(n6187), .O(n6188));
  andx  g05554(.a(n5895), .b(n5738), .O(n6189));
  andx  g05555(.a(n5889), .b(n5728), .O(n6190));
  orx   g05556(.a(n6190), .b(n6189), .O(n6191));
  invx  g05557(.a(n6179), .O(n6192));
  andx  g05558(.a(n6192), .b(n6164), .O(n6193));
  andx  g05559(.a(n6192), .b(n6173), .O(n6194));
  orx   g05560(.a(n6194), .b(n6193), .O(n6195));
  orx   g05561(.a(n6195), .b(n6174), .O(n6196));
  andx  g05562(.a(n6196), .b(n6191), .O(n6197));
  andx  g05563(.a(n5947), .b(n4114), .O(n6198));
  invx  g05564(.a(n6198), .O(n6199));
  orx   g05565(.a(n6199), .b(n6197), .O(n6200));
  andx  g05566(.a(n6200), .b(n6188), .O(n6201));
  orx   g05567(.a(n6201), .b(n5878), .O(n6202));
  orx   g05568(.a(n5754), .b(n5751), .O(n6203));
  orx   g05569(.a(n5753), .b(n5741), .O(n6204));
  andx  g05570(.a(n6204), .b(n6203), .O(n6205));
  andx  g05571(.a(n6205), .b(n5450), .O(n6206));
  andx  g05572(.a(n5753), .b(n5741), .O(n6207));
  andx  g05573(.a(n5754), .b(n5751), .O(n6208));
  orx   g05574(.a(n6208), .b(n6207), .O(n6209));
  andx  g05575(.a(n6209), .b(n5746), .O(n6210));
  orx   g05576(.a(n6210), .b(n6206), .O(n6211));
  andx  g05577(.a(n5947), .b(n4490), .O(n6212));
  invx  g05578(.a(n6212), .O(n6213));
  andx  g05579(.a(n6213), .b(n6201), .O(n6214));
  orx   g05580(.a(n6214), .b(n6211), .O(n6215));
  andx  g05581(.a(n6215), .b(n6202), .O(n6216));
  orx   g05582(.a(n6186), .b(n5897), .O(n6218));
  andx  g05583(.a(n6198), .b(n6218), .O(n6219));
  orx   g05584(.a(n6219), .b(n6187), .O(n6220));
  andx  g05585(.a(n6220), .b(n4490), .O(n6221));
  orx   g05586(.a(n6209), .b(n5746), .O(n6222));
  orx   g05587(.a(n6205), .b(n5450), .O(n6223));
  andx  g05588(.a(n6223), .b(n6222), .O(n6224));
  orx   g05589(.a(n6212), .b(n6220), .O(n6225));
  andx  g05590(.a(n6225), .b(n6224), .O(n6226));
  orx   g05591(.a(n6226), .b(n6221), .O(n6227));
  andx  g05592(.a(n5947), .b(n2724), .O(n6228));
  orx   g05593(.a(n6228), .b(n6227), .O(n6229));
  orx   g05594(.a(n6229), .b(n5876), .O(n6231));
  orx   g05595(.a(n5874), .b(n5763), .O(n6232));
  orx   g05596(.a(n5870), .b(n5426), .O(n6233));
  andx  g05597(.a(n6233), .b(n6232), .O(n6234));
  invx  g05598(.a(n6228), .O(n6236));
  andx  g05599(.a(n6236), .b(n6216), .O(n6237));
  orx   g05600(.a(n6237), .b(n6234), .O(n6239));
  andx  g05601(.a(n6239), .b(n6231), .O(n6240));
  andx  g05602(.a(n6225), .b(n6202), .O(n6241));
  orx   g05603(.a(n6241), .b(n6224), .O(n6242));
  orx   g05604(.a(n6214), .b(n6221), .O(n6243));
  orx   g05605(.a(n6243), .b(n6211), .O(n6244));
  andx  g05606(.a(n6244), .b(n6242), .O(n6245));
  andx  g05607(.a(n148), .b(pi02), .O(n6246));
  andx  g05608(.a(n67), .b(pi00), .O(n6247));
  andx  g05609(.a(n153), .b(pi03), .O(n6248));
  orx   g05610(.a(n6248), .b(n6247), .O(n6249));
  orx   g05611(.a(n6249), .b(n6246), .O(n6250));
  andx  g05612(.a(n159), .b(pi01), .O(n6251));
  andx  g05613(.a(n161), .b(pi05), .O(n6252));
  andx  g05614(.a(n165), .b(pi04), .O(n6253));
  andx  g05615(.a(pi19), .b(pi07), .O(n6254));
  andx  g05616(.a(n103), .b(pi06), .O(n6255));
  orx   g05617(.a(n6255), .b(n6254), .O(n6256));
  orx   g05618(.a(n6256), .b(n6253), .O(n6257));
  orx   g05619(.a(n6257), .b(n6252), .O(n6258));
  orx   g05620(.a(n6258), .b(n6251), .O(n6259));
  orx   g05621(.a(n6259), .b(n6250), .O(n6260));
  andx  g05622(.a(n6260), .b(n92), .O(n6261));
  andx  g05623(.a(n6261), .b(n2724), .O(n6262));
  orx   g05624(.a(n6192), .b(n6164), .O(n6273));
  andx  g05625(.a(n6273), .b(n6180), .O(n6274));
  andx  g05626(.a(n6274), .b(n6183), .O(n6275));
  andx  g05627(.a(n6179), .b(n6178), .O(n6279));
  orx   g05628(.a(n6279), .b(n6193), .O(n6280));
  andx  g05629(.a(n6280), .b(n6173), .O(n6281));
  orx   g05630(.a(n6281), .b(n6275), .O(n6282));
  andx  g05631(.a(n6100), .b(n6099), .O(n6292));
  orx   g05632(.a(n6292), .b(n6116), .O(n6293));
  orx   g05633(.a(n6293), .b(n6094), .O(n6294));
  orx   g05634(.a(n6115), .b(n6085), .O(n6298));
  andx  g05635(.a(n6298), .b(n6101), .O(n6299));
  orx   g05636(.a(n6299), .b(n6104), .O(n6300));
  andx  g05637(.a(n6300), .b(n6294), .O(n6301));
  andx  g05638(.a(n6057), .b(n6035), .O(n6302));
  andx  g05639(.a(n6056), .b(n6079), .O(n6303));
  orx   g05640(.a(n6303), .b(n6302), .O(n6304));
  orx   g05641(.a(n6304), .b(n6054), .O(n6305));
  orx   g05642(.a(n6056), .b(n6079), .O(n6306));
  orx   g05643(.a(n6057), .b(n6035), .O(n6307));
  andx  g05644(.a(n6307), .b(n6306), .O(n6308));
  orx   g05645(.a(n6308), .b(n6082), .O(n6309));
  andx  g05646(.a(n6309), .b(n6305), .O(n6310));
  andx  g05647(.a(n6072), .b(n6071), .O(n6320));
  orx   g05648(.a(n6320), .b(n6032), .O(n6321));
  orx   g05649(.a(n6321), .b(n6029), .O(n6322));
  orx   g05650(.a(n6031), .b(n6020), .O(n6326));
  andx  g05651(.a(n6326), .b(n6073), .O(n6327));
  orx   g05652(.a(n6327), .b(n6076), .O(n6328));
  andx  g05653(.a(n6328), .b(n6322), .O(n6329));
  orx   g05654(.a(n6068), .b(n6006), .O(n6330));
  orx   g05655(.a(n6017), .b(n6063), .O(n6331));
  andx  g05656(.a(n6331), .b(n6330), .O(n6332));
  orx   g05657(.a(n6332), .b(n6015), .O(n6333));
  andx  g05658(.a(n6017), .b(n6063), .O(n6334));
  andx  g05659(.a(n6068), .b(n6006), .O(n6335));
  orx   g05660(.a(n6335), .b(n6334), .O(n6336));
  orx   g05661(.a(n6336), .b(n6066), .O(n6337));
  andx  g05662(.a(n6337), .b(n6333), .O(n6338));
  andx  g05663(.a(n6004), .b(n5982), .O(n6339));
  andx  g05664(.a(n6061), .b(n6001), .O(n6340));
  orx   g05665(.a(n6340), .b(n6339), .O(n6341));
  andx  g05666(.a(n6341), .b(n5987), .O(n6342));
  orx   g05667(.a(n6061), .b(n6001), .O(n6343));
  orx   g05668(.a(n6004), .b(n5982), .O(n6344));
  andx  g05669(.a(n6344), .b(n6343), .O(n6345));
  andx  g05670(.a(n6345), .b(n5924), .O(n6346));
  orx   g05671(.a(n6346), .b(n6342), .O(n6347));
  orx   g05672(.a(n5979), .b(n5998), .O(n6348));
  orx   g05673(.a(n5989), .b(n5977), .O(n6349));
  andx  g05674(.a(n6349), .b(n6348), .O(n6350));
  orx   g05675(.a(n6350), .b(n5992), .O(n6351));
  andx  g05676(.a(n5989), .b(n5977), .O(n6352));
  andx  g05677(.a(n5979), .b(n5998), .O(n6353));
  orx   g05678(.a(n6353), .b(n6352), .O(n6354));
  orx   g05679(.a(n6354), .b(n5929), .O(n6355));
  andx  g05680(.a(n6355), .b(n6351), .O(n6356));
  orx   g05681(.a(n5996), .b(n5962), .O(n6357));
  andx  g05682(.a(n6357), .b(n5973), .O(n6358));
  andx  g05683(.a(n5975), .b(n5993), .O(n6359));
  andx  g05684(.a(n6359), .b(n5995), .O(n6360));
  orx   g05685(.a(n6360), .b(n6358), .O(n6361));
  andx  g05686(.a(n6261), .b(n3230), .O(n6362));
  invx  g05687(.a(n5956), .O(n6363));
  andx  g05688(.a(n6363), .b(n5955), .O(n6364));
  invx  g05689(.a(n5955), .O(n6365));
  andx  g05690(.a(n5956), .b(n6365), .O(n6366));
  orx   g05691(.a(n6366), .b(n6364), .O(n6367));
  andx  g05692(.a(n6367), .b(n6362), .O(n6368));
  andx  g05693(.a(n5947), .b(n1790), .O(n6369));
  andx  g05694(.a(n6261), .b(n3258), .O(n6370));
  andx  g05695(.a(n6370), .b(n6369), .O(n6371));
  andx  g05696(.a(n6371), .b(n6362), .O(n6372));
  andx  g05697(.a(n6371), .b(n6367), .O(n6373));
  orx   g05698(.a(n6373), .b(n6372), .O(n6374));
  orx   g05699(.a(n6374), .b(n6368), .O(n6375));
  andx  g05700(.a(n6375), .b(n3221), .O(n6376));
  invx  g05701(.a(n5957), .O(n6377));
  andx  g05702(.a(n6377), .b(n5948), .O(n6378));
  invx  g05703(.a(n6378), .O(n6379));
  orx   g05704(.a(n6377), .b(n5948), .O(n6380));
  andx  g05705(.a(n6380), .b(n6379), .O(n6381));
  andx  g05706(.a(n5949), .b(n5951), .O(n6382));
  orx   g05707(.a(n6382), .b(n5566), .O(n6383));
  andx  g05708(.a(n6383), .b(n6381), .O(n6384));
  invx  g05709(.a(n6384), .O(n6385));
  orx   g05710(.a(n6383), .b(n6381), .O(n6386));
  andx  g05711(.a(n6386), .b(n6385), .O(n6387));
  andx  g05712(.a(n6261), .b(n3221), .O(n6388));
  orx   g05713(.a(n6388), .b(n6375), .O(n6389));
  andx  g05714(.a(n6389), .b(n6387), .O(n6390));
  orx   g05715(.a(n6390), .b(n6376), .O(n6391));
  andx  g05716(.a(n6391), .b(n6361), .O(n6392));
  andx  g05717(.a(n6261), .b(n3210), .O(n6393));
  orx   g05718(.a(n6391), .b(n6361), .O(n6394));
  andx  g05719(.a(n6394), .b(n6393), .O(n6395));
  orx   g05720(.a(n6395), .b(n6392), .O(n6396));
  andx  g05721(.a(n6396), .b(n6356), .O(n6397));
  orx   g05722(.a(n6396), .b(n6356), .O(n6398));
  andx  g05723(.a(n6261), .b(n3284), .O(n6399));
  andx  g05724(.a(n6399), .b(n6398), .O(n6400));
  orx   g05725(.a(n6400), .b(n6397), .O(n6401));
  andx  g05726(.a(n6401), .b(n6347), .O(n6402));
  andx  g05727(.a(n6261), .b(n3180), .O(n6403));
  orx   g05728(.a(n6401), .b(n6347), .O(n6404));
  andx  g05729(.a(n6404), .b(n6403), .O(n6405));
  orx   g05730(.a(n6405), .b(n6402), .O(n6406));
  andx  g05731(.a(n6406), .b(n6338), .O(n6407));
  orx   g05732(.a(n6406), .b(n6338), .O(n6408));
  andx  g05733(.a(n6261), .b(n3429), .O(n6409));
  andx  g05734(.a(n6409), .b(n6408), .O(n6410));
  orx   g05735(.a(n6410), .b(n6407), .O(n6411));
  andx  g05736(.a(n6411), .b(n6329), .O(n6412));
  andx  g05737(.a(n6261), .b(n3171), .O(n6413));
  orx   g05738(.a(n6411), .b(n6329), .O(n6414));
  andx  g05739(.a(n6414), .b(n6413), .O(n6415));
  orx   g05740(.a(n6415), .b(n6412), .O(n6416));
  andx  g05741(.a(n6416), .b(n6310), .O(n6417));
  orx   g05742(.a(n6416), .b(n6310), .O(n6418));
  andx  g05743(.a(n6261), .b(n3413), .O(n6419));
  andx  g05744(.a(n6419), .b(n6418), .O(n6420));
  orx   g05745(.a(n6420), .b(n6417), .O(n6421));
  andx  g05746(.a(n6421), .b(n6301), .O(n6422));
  invx  g05747(.a(n6422), .O(n6423));
  andx  g05748(.a(n6261), .b(n3645), .O(n6424));
  invx  g05749(.a(n6424), .O(n6425));
  andx  g05750(.a(n6299), .b(n6104), .O(n6426));
  andx  g05751(.a(n6293), .b(n6094), .O(n6427));
  orx   g05752(.a(n6427), .b(n6426), .O(n6428));
  invx  g05753(.a(n6417), .O(n6429));
  andx  g05754(.a(n6308), .b(n6082), .O(n6430));
  andx  g05755(.a(n6304), .b(n6054), .O(n6431));
  orx   g05756(.a(n6431), .b(n6430), .O(n6432));
  andx  g05757(.a(n6327), .b(n6076), .O(n6433));
  andx  g05758(.a(n6321), .b(n6029), .O(n6434));
  orx   g05759(.a(n6434), .b(n6433), .O(n6435));
  invx  g05760(.a(n6407), .O(n6436));
  andx  g05761(.a(n6336), .b(n6066), .O(n6437));
  andx  g05762(.a(n6332), .b(n6015), .O(n6438));
  orx   g05763(.a(n6438), .b(n6437), .O(n6439));
  invx  g05764(.a(n6402), .O(n6440));
  invx  g05765(.a(n6403), .O(n6441));
  orx   g05766(.a(n6345), .b(n5924), .O(n6442));
  orx   g05767(.a(n6341), .b(n5987), .O(n6443));
  andx  g05768(.a(n6443), .b(n6442), .O(n6444));
  invx  g05769(.a(n6397), .O(n6445));
  andx  g05770(.a(n6354), .b(n5929), .O(n6446));
  andx  g05771(.a(n6350), .b(n5992), .O(n6447));
  orx   g05772(.a(n6447), .b(n6446), .O(n6448));
  invx  g05773(.a(n6392), .O(n6449));
  invx  g05774(.a(n6393), .O(n6450));
  orx   g05775(.a(n6359), .b(n5995), .O(n6451));
  orx   g05776(.a(n6357), .b(n5973), .O(n6452));
  andx  g05777(.a(n6452), .b(n6451), .O(n6453));
  invx  g05778(.a(n6376), .O(n6454));
  invx  g05779(.a(n6386), .O(n6455));
  orx   g05780(.a(n6455), .b(n6384), .O(n6456));
  invx  g05781(.a(n6389), .O(n6457));
  orx   g05782(.a(n6457), .b(n6456), .O(n6458));
  andx  g05783(.a(n6458), .b(n6454), .O(n6459));
  andx  g05784(.a(n6459), .b(n6453), .O(n6460));
  orx   g05785(.a(n6460), .b(n6450), .O(n6461));
  andx  g05786(.a(n6461), .b(n6449), .O(n6462));
  andx  g05787(.a(n6462), .b(n6448), .O(n6463));
  invx  g05788(.a(n6399), .O(n6464));
  orx   g05789(.a(n6464), .b(n6463), .O(n6465));
  andx  g05790(.a(n6465), .b(n6445), .O(n6466));
  andx  g05791(.a(n6466), .b(n6444), .O(n6467));
  orx   g05792(.a(n6467), .b(n6441), .O(n6468));
  andx  g05793(.a(n6468), .b(n6440), .O(n6469));
  andx  g05794(.a(n6469), .b(n6439), .O(n6470));
  invx  g05795(.a(n6409), .O(n6471));
  orx   g05796(.a(n6471), .b(n6470), .O(n6472));
  andx  g05797(.a(n6472), .b(n6436), .O(n6473));
  orx   g05798(.a(n6473), .b(n6435), .O(n6474));
  invx  g05799(.a(n6261), .O(n6475));
  orx   g05800(.a(n6475), .b(n3418), .O(n6476));
  andx  g05801(.a(n6473), .b(n6435), .O(n6477));
  orx   g05802(.a(n6477), .b(n6476), .O(n6478));
  andx  g05803(.a(n6478), .b(n6474), .O(n6479));
  andx  g05804(.a(n6479), .b(n6432), .O(n6480));
  orx   g05805(.a(n6475), .b(n4989), .O(n6481));
  orx   g05806(.a(n6481), .b(n6480), .O(n6482));
  andx  g05807(.a(n6482), .b(n6429), .O(n6483));
  andx  g05808(.a(n6483), .b(n6428), .O(n6484));
  orx   g05809(.a(n6484), .b(n6425), .O(n6485));
  andx  g05810(.a(n6485), .b(n6423), .O(n6486));
  andx  g05811(.a(n6111), .b(n6119), .O(n6487));
  andx  g05812(.a(n6110), .b(n6107), .O(n6488));
  orx   g05813(.a(n6488), .b(n6487), .O(n6489));
  orx   g05814(.a(n6489), .b(n5915), .O(n6490));
  orx   g05815(.a(n6110), .b(n6107), .O(n6491));
  orx   g05816(.a(n6111), .b(n6119), .O(n6492));
  andx  g05817(.a(n6492), .b(n6491), .O(n6493));
  orx   g05818(.a(n6493), .b(n6114), .O(n6494));
  andx  g05819(.a(n6494), .b(n6490), .O(n6495));
  andx  g05820(.a(n6495), .b(n6486), .O(n6496));
  andx  g05821(.a(n6261), .b(n3721), .O(n6497));
  invx  g05822(.a(n6497), .O(n6498));
  orx   g05823(.a(n6498), .b(n6496), .O(n6499));
  orx   g05824(.a(n6421), .b(n6301), .O(n6500));
  andx  g05825(.a(n6500), .b(n6424), .O(n6501));
  orx   g05826(.a(n6501), .b(n6422), .O(n6502));
  andx  g05827(.a(n6493), .b(n6114), .O(n6503));
  andx  g05828(.a(n6489), .b(n5915), .O(n6504));
  orx   g05829(.a(n6504), .b(n6503), .O(n6505));
  andx  g05830(.a(n6505), .b(n6502), .O(n6506));
  invx  g05831(.a(n6506), .O(n6507));
  andx  g05832(.a(n6507), .b(n6499), .O(n6508));
  andx  g05833(.a(n6153), .b(n6158), .O(n6509));
  andx  g05834(.a(n6154), .b(n6122), .O(n6510));
  orx   g05835(.a(n6510), .b(n6509), .O(n6511));
  andx  g05836(.a(n6511), .b(n6151), .O(n6512));
  orx   g05837(.a(n6154), .b(n6122), .O(n6513));
  orx   g05838(.a(n6153), .b(n6158), .O(n6514));
  andx  g05839(.a(n6514), .b(n6513), .O(n6515));
  andx  g05840(.a(n6515), .b(n6161), .O(n6516));
  orx   g05841(.a(n6516), .b(n6512), .O(n6517));
  andx  g05842(.a(n6517), .b(n6508), .O(n6518));
  andx  g05843(.a(n6261), .b(n4063), .O(n6519));
  invx  g05844(.a(n6519), .O(n6520));
  andx  g05845(.a(n6520), .b(n6508), .O(n6521));
  andx  g05846(.a(n6520), .b(n6517), .O(n6522));
  orx   g05847(.a(n6522), .b(n6521), .O(n6523));
  orx   g05848(.a(n6523), .b(n6518), .O(n6524));
  andx  g05849(.a(n6524), .b(n6282), .O(n6525));
  andx  g05850(.a(n6261), .b(n4114), .O(n6526));
  invx  g05851(.a(n6526), .O(n6527));
  orx   g05852(.a(n6527), .b(n6525), .O(n6528));
  orx   g05853(.a(n6280), .b(n6173), .O(n6529));
  orx   g05854(.a(n6274), .b(n6183), .O(n6530));
  andx  g05855(.a(n6530), .b(n6529), .O(n6531));
  invx  g05856(.a(n6518), .O(n6532));
  orx   g05857(.a(n6505), .b(n6502), .O(n6533));
  andx  g05858(.a(n6497), .b(n6533), .O(n6534));
  orx   g05859(.a(n6506), .b(n6534), .O(n6535));
  orx   g05860(.a(n6519), .b(n6535), .O(n6536));
  orx   g05861(.a(n6515), .b(n6161), .O(n6537));
  orx   g05862(.a(n6511), .b(n6151), .O(n6538));
  andx  g05863(.a(n6538), .b(n6537), .O(n6539));
  orx   g05864(.a(n6519), .b(n6539), .O(n6540));
  andx  g05865(.a(n6540), .b(n6536), .O(n6541));
  andx  g05866(.a(n6541), .b(n6532), .O(n6542));
  andx  g05867(.a(n6542), .b(n6531), .O(n6543));
  invx  g05868(.a(n6543), .O(n6544));
  andx  g05869(.a(n6544), .b(n6528), .O(n6545));
  andx  g05870(.a(n6199), .b(n6186), .O(n6546));
  andx  g05871(.a(n6198), .b(n6196), .O(n6547));
  orx   g05872(.a(n6547), .b(n6546), .O(n6548));
  orx   g05873(.a(n6548), .b(n6191), .O(n6549));
  orx   g05874(.a(n6198), .b(n6196), .O(n6550));
  orx   g05875(.a(n6199), .b(n6186), .O(n6551));
  andx  g05876(.a(n6551), .b(n6550), .O(n6552));
  orx   g05877(.a(n6552), .b(n5897), .O(n6553));
  andx  g05878(.a(n6553), .b(n6549), .O(n6554));
  andx  g05879(.a(n6554), .b(n6545), .O(n6555));
  invx  g05880(.a(n6555), .O(n6556));
  orx   g05881(.a(n6542), .b(n6531), .O(n6557));
  andx  g05882(.a(n6526), .b(n6557), .O(n6558));
  orx   g05883(.a(n6543), .b(n6558), .O(n6559));
  andx  g05884(.a(n6261), .b(n4490), .O(n6560));
  orx   g05885(.a(n6560), .b(n6559), .O(n6561));
  andx  g05886(.a(n6552), .b(n5897), .O(n6562));
  andx  g05887(.a(n6548), .b(n6191), .O(n6563));
  orx   g05888(.a(n6563), .b(n6562), .O(n6564));
  orx   g05889(.a(n6560), .b(n6564), .O(n6565));
  andx  g05890(.a(n6565), .b(n6561), .O(n6566));
  andx  g05891(.a(n6566), .b(n6556), .O(n6567));
  andx  g05892(.a(n6567), .b(n6245), .O(n6568));
  andx  g05893(.a(n6568), .b(n6240), .O(n6572));
  andx  g05894(.a(n6229), .b(n5876), .O(n6573));
  andx  g05895(.a(n5414), .b(n5413), .O(n6576));
  andx  g05896(.a(n5409), .b(n5364), .O(n6577));
  orx   g05897(.a(n6577), .b(n6576), .O(n6578));
  orx   g05898(.a(n5772), .b(n5769), .O(n6579));
  invx  g05899(.a(n6579), .O(n6580));
  orx   g05900(.a(n5772), .b(n6580), .O(n6582));
  andx  g05901(.a(n6582), .b(n6578), .O(n6583));
  invx  g05902(.a(n5772), .O(n6584));
  andx  g05903(.a(n6584), .b(n6579), .O(n6585));
  andx  g05904(.a(n6585), .b(n5416), .O(n6586));
  orx   g05905(.a(n6586), .b(n6583), .O(n6587));
  andx  g05906(.a(n6587), .b(n6239), .O(n6588));
  orx   g05907(.a(n6585), .b(n5416), .O(n6589));
  orx   g05908(.a(n6582), .b(n6578), .O(n6590));
  andx  g05909(.a(n6590), .b(n6589), .O(n6591));
  andx  g05910(.a(n6591), .b(n6573), .O(n6592));
  orx   g05911(.a(n6592), .b(n6588), .O(n6593));
  orx   g05912(.a(n6593), .b(n6572), .O(n6594));
  andx  g05913(.a(n159), .b(pi00), .O(n6595));
  andx  g05914(.a(n165), .b(pi03), .O(n6596));
  andx  g05915(.a(n161), .b(pi04), .O(n6597));
  andx  g05916(.a(n103), .b(pi05), .O(n6598));
  andx  g05917(.a(pi19), .b(pi06), .O(n6599));
  orx   g05918(.a(n6599), .b(n6598), .O(n6600));
  orx   g05919(.a(n6600), .b(n6597), .O(n6601));
  orx   g05920(.a(n6601), .b(n6596), .O(n6602));
  andx  g05921(.a(n148), .b(pi01), .O(n6603));
  andx  g05922(.a(n153), .b(pi02), .O(n6604));
  orx   g05923(.a(n6604), .b(n6603), .O(n6605));
  orx   g05924(.a(n6605), .b(n6602), .O(n6606));
  orx   g05925(.a(n6606), .b(n6595), .O(n6607));
  andx  g05926(.a(n6607), .b(n2724), .O(n6608));
  invx  g05927(.a(n6608), .O(n6609));
  invx  g05928(.a(n6560), .O(n6619));
  orx   g05929(.a(n6619), .b(n6545), .O(n6620));
  andx  g05930(.a(n6620), .b(n6561), .O(n6621));
  andx  g05931(.a(n6621), .b(n6564), .O(n6622));
  andx  g05932(.a(n6619), .b(n6545), .O(n6626));
  andx  g05933(.a(n6560), .b(n6559), .O(n6627));
  orx   g05934(.a(n6627), .b(n6626), .O(n6628));
  andx  g05935(.a(n6628), .b(n6554), .O(n6629));
  orx   g05936(.a(n6629), .b(n6622), .O(n6630));
  orx   g05937(.a(n6497), .b(n6486), .O(n6631));
  orx   g05938(.a(n6498), .b(n6502), .O(n6632));
  andx  g05939(.a(n6632), .b(n6631), .O(n6633));
  orx   g05940(.a(n6633), .b(n6495), .O(n6634));
  andx  g05941(.a(n6498), .b(n6502), .O(n6635));
  andx  g05942(.a(n6497), .b(n6486), .O(n6636));
  orx   g05943(.a(n6636), .b(n6635), .O(n6637));
  orx   g05944(.a(n6637), .b(n6505), .O(n6638));
  andx  g05945(.a(n6638), .b(n6634), .O(n6639));
  orx   g05946(.a(n6424), .b(n6483), .O(n6640));
  orx   g05947(.a(n6425), .b(n6421), .O(n6641));
  andx  g05948(.a(n6641), .b(n6640), .O(n6642));
  andx  g05949(.a(n6642), .b(n6428), .O(n6643));
  andx  g05950(.a(n6425), .b(n6421), .O(n6644));
  andx  g05951(.a(n6424), .b(n6483), .O(n6645));
  orx   g05952(.a(n6645), .b(n6644), .O(n6646));
  andx  g05953(.a(n6646), .b(n6301), .O(n6647));
  orx   g05954(.a(n6647), .b(n6643), .O(n6648));
  orx   g05955(.a(n6419), .b(n6479), .O(n6649));
  orx   g05956(.a(n6481), .b(n6416), .O(n6650));
  andx  g05957(.a(n6650), .b(n6649), .O(n6651));
  orx   g05958(.a(n6651), .b(n6310), .O(n6652));
  andx  g05959(.a(n6481), .b(n6416), .O(n6653));
  andx  g05960(.a(n6419), .b(n6479), .O(n6654));
  orx   g05961(.a(n6654), .b(n6653), .O(n6655));
  orx   g05962(.a(n6655), .b(n6432), .O(n6656));
  andx  g05963(.a(n6656), .b(n6652), .O(n6657));
  andx  g05964(.a(n6476), .b(n6411), .O(n6658));
  andx  g05965(.a(n6413), .b(n6473), .O(n6659));
  orx   g05966(.a(n6659), .b(n6658), .O(n6660));
  orx   g05967(.a(n6660), .b(n6435), .O(n6661));
  orx   g05968(.a(n6413), .b(n6473), .O(n6662));
  orx   g05969(.a(n6476), .b(n6411), .O(n6663));
  andx  g05970(.a(n6663), .b(n6662), .O(n6664));
  orx   g05971(.a(n6664), .b(n6329), .O(n6665));
  andx  g05972(.a(n6665), .b(n6661), .O(n6666));
  orx   g05973(.a(n6409), .b(n6469), .O(n6667));
  orx   g05974(.a(n6471), .b(n6406), .O(n6668));
  andx  g05975(.a(n6668), .b(n6667), .O(n6669));
  orx   g05976(.a(n6669), .b(n6338), .O(n6670));
  andx  g05977(.a(n6471), .b(n6406), .O(n6671));
  andx  g05978(.a(n6409), .b(n6469), .O(n6672));
  orx   g05979(.a(n6672), .b(n6671), .O(n6673));
  orx   g05980(.a(n6673), .b(n6439), .O(n6674));
  andx  g05981(.a(n6674), .b(n6670), .O(n6675));
  orx   g05982(.a(n6399), .b(n6462), .O(n6676));
  orx   g05983(.a(n6464), .b(n6396), .O(n6677));
  andx  g05984(.a(n6677), .b(n6676), .O(n6678));
  orx   g05985(.a(n6678), .b(n6356), .O(n6679));
  andx  g05986(.a(n6464), .b(n6396), .O(n6680));
  andx  g05987(.a(n6399), .b(n6462), .O(n6681));
  orx   g05988(.a(n6681), .b(n6680), .O(n6682));
  orx   g05989(.a(n6682), .b(n6448), .O(n6683));
  andx  g05990(.a(n6683), .b(n6679), .O(n6684));
  andx  g05991(.a(n6450), .b(n6391), .O(n6685));
  andx  g05992(.a(n6393), .b(n6459), .O(n6686));
  orx   g05993(.a(n6686), .b(n6685), .O(n6687));
  andx  g05994(.a(n6687), .b(n6453), .O(n6688));
  orx   g05995(.a(n6393), .b(n6459), .O(n6689));
  orx   g05996(.a(n6450), .b(n6391), .O(n6690));
  andx  g05997(.a(n6690), .b(n6689), .O(n6691));
  andx  g05998(.a(n6691), .b(n6361), .O(n6692));
  orx   g05999(.a(n6692), .b(n6688), .O(n6693));
  andx  g06000(.a(n6389), .b(n6454), .O(n6694));
  orx   g06001(.a(n6694), .b(n6456), .O(n6695));
  invx  g06002(.a(n6695), .O(n6696));
  andx  g06003(.a(n6694), .b(n6456), .O(n6697));
  orx   g06004(.a(n6697), .b(n6696), .O(n6698));
  andx  g06005(.a(n6607), .b(n3230), .O(n6699));
  invx  g06006(.a(n6369), .O(n6700));
  orx   g06007(.a(n6370), .b(n6700), .O(n6701));
  andx  g06008(.a(n6370), .b(n6700), .O(n6702));
  invx  g06009(.a(n6702), .O(n6703));
  andx  g06010(.a(n6703), .b(n6701), .O(n6704));
  andx  g06011(.a(n7028), .b(n6699), .O(n6706));
  andx  g06012(.a(n6607), .b(n3258), .O(n6707));
  andx  g06013(.a(n6261), .b(n1790), .O(n6708));
  andx  g06014(.a(n6708), .b(n6707), .O(n6709));
  andx  g06015(.a(n6709), .b(n6699), .O(n6710));
  andx  g06016(.a(n6709), .b(n7028), .O(n6711));
  orx   g06017(.a(n6711), .b(n6710), .O(n6712));
  orx   g06018(.a(n6712), .b(n6706), .O(n6713));
  andx  g06019(.a(n6713), .b(n3221), .O(n6714));
  andx  g06020(.a(n6363), .b(n6365), .O(n6715));
  orx   g06021(.a(n6715), .b(n5957), .O(n6716));
  invx  g06022(.a(n6372), .O(n6717));
  orx   g06023(.a(n6371), .b(n6362), .O(n6718));
  andx  g06024(.a(n6718), .b(n6717), .O(n6719));
  invx  g06025(.a(n6719), .O(n6720));
  andx  g06026(.a(n6720), .b(n6716), .O(n6721));
  invx  g06027(.a(n6721), .O(n6722));
  orx   g06028(.a(n6720), .b(n6716), .O(n6723));
  andx  g06029(.a(n6723), .b(n6722), .O(n6724));
  andx  g06030(.a(n6607), .b(n3221), .O(n6725));
  orx   g06031(.a(n6725), .b(n6713), .O(n6726));
  andx  g06032(.a(n6726), .b(n6724), .O(n6727));
  orx   g06033(.a(n6727), .b(n6714), .O(n6728));
  andx  g06034(.a(n6728), .b(n6698), .O(n6729));
  andx  g06035(.a(n6607), .b(n3210), .O(n6730));
  orx   g06036(.a(n6728), .b(n6698), .O(n6731));
  andx  g06037(.a(n6731), .b(n6730), .O(n6732));
  orx   g06038(.a(n6732), .b(n6729), .O(n6733));
  andx  g06039(.a(n6733), .b(n6693), .O(n6734));
  invx  g06040(.a(n6734), .O(n6735));
  orx   g06041(.a(n6691), .b(n6361), .O(n6736));
  orx   g06042(.a(n6687), .b(n6453), .O(n6737));
  andx  g06043(.a(n6737), .b(n6736), .O(n6738));
  invx  g06044(.a(n6729), .O(n6739));
  invx  g06045(.a(n6730), .O(n6740));
  invx  g06046(.a(n6697), .O(n6741));
  andx  g06047(.a(n6741), .b(n6695), .O(n6742));
  invx  g06048(.a(n6714), .O(n6743));
  invx  g06049(.a(n6723), .O(n6744));
  orx   g06050(.a(n6744), .b(n6721), .O(n6745));
  invx  g06051(.a(n6726), .O(n6746));
  orx   g06052(.a(n6746), .b(n6745), .O(n6747));
  andx  g06053(.a(n6747), .b(n6743), .O(n6748));
  andx  g06054(.a(n6748), .b(n6742), .O(n6749));
  orx   g06055(.a(n6749), .b(n6740), .O(n6750));
  andx  g06056(.a(n6750), .b(n6739), .O(n6751));
  andx  g06057(.a(n6751), .b(n6738), .O(n6752));
  andx  g06058(.a(n6607), .b(n3284), .O(n6753));
  invx  g06059(.a(n6753), .O(n6754));
  orx   g06060(.a(n6754), .b(n6752), .O(n6755));
  andx  g06061(.a(n6755), .b(n6735), .O(n6756));
  andx  g06062(.a(n6756), .b(n6684), .O(n6757));
  andx  g06063(.a(n6607), .b(n3180), .O(n6758));
  invx  g06064(.a(n6758), .O(n6759));
  orx   g06065(.a(n6759), .b(n6757), .O(n6760));
  andx  g06066(.a(n6682), .b(n6448), .O(n6761));
  andx  g06067(.a(n6678), .b(n6356), .O(n6762));
  orx   g06068(.a(n6762), .b(n6761), .O(n6763));
  orx   g06069(.a(n6733), .b(n6693), .O(n6764));
  andx  g06070(.a(n6753), .b(n6764), .O(n6765));
  orx   g06071(.a(n6765), .b(n6734), .O(n6766));
  andx  g06072(.a(n6766), .b(n6763), .O(n6767));
  invx  g06073(.a(n6767), .O(n6768));
  andx  g06074(.a(n6768), .b(n6760), .O(n6769));
  orx   g06075(.a(n6403), .b(n6466), .O(n6770));
  orx   g06076(.a(n6441), .b(n6401), .O(n6771));
  andx  g06077(.a(n6771), .b(n6770), .O(n6772));
  andx  g06078(.a(n6772), .b(n6444), .O(n6773));
  andx  g06079(.a(n6441), .b(n6401), .O(n6774));
  andx  g06080(.a(n6403), .b(n6466), .O(n6775));
  orx   g06081(.a(n6775), .b(n6774), .O(n6776));
  andx  g06082(.a(n6776), .b(n6347), .O(n6777));
  orx   g06083(.a(n6777), .b(n6773), .O(n6778));
  andx  g06084(.a(n6778), .b(n6769), .O(n6779));
  andx  g06085(.a(n6607), .b(n3429), .O(n6780));
  invx  g06086(.a(n6780), .O(n6781));
  andx  g06087(.a(n6781), .b(n6769), .O(n6782));
  andx  g06088(.a(n6781), .b(n6778), .O(n6783));
  orx   g06089(.a(n6783), .b(n6782), .O(n6784));
  orx   g06090(.a(n6784), .b(n6779), .O(n6785));
  andx  g06091(.a(n6785), .b(n6675), .O(n6786));
  andx  g06092(.a(n6607), .b(n3171), .O(n6787));
  invx  g06093(.a(n6787), .O(n6788));
  orx   g06094(.a(n6788), .b(n6786), .O(n6789));
  andx  g06095(.a(n6673), .b(n6439), .O(n6790));
  andx  g06096(.a(n6669), .b(n6338), .O(n6791));
  orx   g06097(.a(n6791), .b(n6790), .O(n6792));
  invx  g06098(.a(n6779), .O(n6793));
  orx   g06099(.a(n6766), .b(n6763), .O(n6794));
  andx  g06100(.a(n6758), .b(n6794), .O(n6795));
  orx   g06101(.a(n6767), .b(n6795), .O(n6796));
  orx   g06102(.a(n6780), .b(n6796), .O(n6797));
  orx   g06103(.a(n6776), .b(n6347), .O(n6798));
  orx   g06104(.a(n6772), .b(n6444), .O(n6799));
  andx  g06105(.a(n6799), .b(n6798), .O(n6800));
  orx   g06106(.a(n6780), .b(n6800), .O(n6801));
  andx  g06107(.a(n6801), .b(n6797), .O(n6802));
  andx  g06108(.a(n6802), .b(n6793), .O(n6803));
  andx  g06109(.a(n6803), .b(n6792), .O(n6804));
  invx  g06110(.a(n6804), .O(n6805));
  andx  g06111(.a(n6805), .b(n6789), .O(n6806));
  andx  g06112(.a(n6806), .b(n6666), .O(n6807));
  andx  g06113(.a(n6607), .b(n3413), .O(n6808));
  invx  g06114(.a(n6808), .O(n6809));
  andx  g06115(.a(n6809), .b(n6666), .O(n6810));
  andx  g06116(.a(n6809), .b(n6806), .O(n6811));
  orx   g06117(.a(n6811), .b(n6810), .O(n6812));
  orx   g06118(.a(n6812), .b(n6807), .O(n6813));
  andx  g06119(.a(n6813), .b(n6657), .O(n6814));
  invx  g06120(.a(n6607), .O(n6815));
  orx   g06121(.a(n6815), .b(n4509), .O(n6816));
  orx   g06122(.a(n6816), .b(n6814), .O(n6817));
  orx   g06123(.a(n6813), .b(n6657), .O(n6818));
  andx  g06124(.a(n6818), .b(n6817), .O(n6819));
  andx  g06125(.a(n6819), .b(n6648), .O(n6820));
  invx  g06126(.a(n6820), .O(n6821));
  orx   g06127(.a(n6646), .b(n6301), .O(n6822));
  orx   g06128(.a(n6642), .b(n6428), .O(n6823));
  andx  g06129(.a(n6823), .b(n6822), .O(n6824));
  andx  g06130(.a(n6607), .b(n3721), .O(n6825));
  orx   g06131(.a(n6825), .b(n6824), .O(n6826));
  orx   g06132(.a(n3719), .b(n3718), .O(n6827));
  orx   g06133(.a(n3714), .b(n3712), .O(n6828));
  andx  g06134(.a(n6828), .b(n6827), .O(n6829));
  orx   g06135(.a(n6815), .b(n6829), .O(n6830));
  andx  g06136(.a(n6830), .b(n6819), .O(n6831));
  invx  g06137(.a(n6831), .O(n6832));
  andx  g06138(.a(n6832), .b(n6826), .O(n6833));
  andx  g06139(.a(n6833), .b(n6821), .O(n6834));
  andx  g06140(.a(n6834), .b(n6639), .O(n6835));
  invx  g06141(.a(n6835), .O(n6836));
  andx  g06142(.a(n6607), .b(n4063), .O(n6837));
  invx  g06143(.a(n6837), .O(n6838));
  andx  g06144(.a(n6637), .b(n6505), .O(n6839));
  andx  g06145(.a(n6633), .b(n6495), .O(n6840));
  orx   g06146(.a(n6840), .b(n6839), .O(n6841));
  andx  g06147(.a(n6830), .b(n6648), .O(n6842));
  orx   g06148(.a(n6831), .b(n6842), .O(n6843));
  orx   g06149(.a(n6843), .b(n6820), .O(n6844));
  andx  g06150(.a(n6844), .b(n6841), .O(n6845));
  orx   g06151(.a(n6845), .b(n6838), .O(n6846));
  andx  g06152(.a(n6846), .b(n6836), .O(n6847));
  orx   g06153(.a(n6520), .b(n6508), .O(n6855));
  andx  g06154(.a(n6855), .b(n6536), .O(n6856));
  andx  g06155(.a(n6856), .b(n6539), .O(n6857));
  andx  g06156(.a(n6519), .b(n6535), .O(n6859));
  orx   g06157(.a(n6859), .b(n6521), .O(n6860));
  andx  g06158(.a(n6860), .b(n6517), .O(n6861));
  orx   g06159(.a(n6861), .b(n6857), .O(n6862));
  andx  g06160(.a(n6862), .b(n6847), .O(n6863));
  andx  g06161(.a(n6607), .b(n4114), .O(n6864));
  invx  g06162(.a(n6864), .O(n6865));
  orx   g06163(.a(n6865), .b(n6863), .O(n6866));
  orx   g06164(.a(n6834), .b(n6639), .O(n6867));
  andx  g06165(.a(n6867), .b(n6837), .O(n6868));
  orx   g06166(.a(n6868), .b(n6835), .O(n6869));
  orx   g06167(.a(n6860), .b(n6517), .O(n6870));
  orx   g06168(.a(n6856), .b(n6539), .O(n6871));
  andx  g06169(.a(n6871), .b(n6870), .O(n6872));
  andx  g06170(.a(n6872), .b(n6869), .O(n6873));
  invx  g06171(.a(n6873), .O(n6874));
  andx  g06172(.a(n6874), .b(n6866), .O(n6875));
  andx  g06173(.a(n6526), .b(n6542), .O(n6876));
  andx  g06174(.a(n6527), .b(n6524), .O(n6877));
  orx   g06175(.a(n6877), .b(n6876), .O(n6878));
  andx  g06176(.a(n6878), .b(n6282), .O(n6879));
  orx   g06177(.a(n6527), .b(n6524), .O(n6880));
  orx   g06178(.a(n6526), .b(n6542), .O(n6881));
  andx  g06179(.a(n6881), .b(n6880), .O(n6882));
  andx  g06180(.a(n6882), .b(n6531), .O(n6883));
  orx   g06181(.a(n6883), .b(n6879), .O(n6884));
  andx  g06182(.a(n6884), .b(n6875), .O(n6885));
  andx  g06183(.a(n6607), .b(n4490), .O(n6886));
  invx  g06184(.a(n6886), .O(n6887));
  andx  g06185(.a(n6887), .b(n6875), .O(n6888));
  andx  g06186(.a(n6887), .b(n6884), .O(n6889));
  orx   g06187(.a(n6889), .b(n6888), .O(n6890));
  orx   g06188(.a(n6890), .b(n6885), .O(n6891));
  orx   g06189(.a(n6628), .b(n6554), .O(n6894));
  orx   g06190(.a(n6621), .b(n6564), .O(n6895));
  andx  g06191(.a(n6895), .b(n6894), .O(n6896));
  invx  g06192(.a(n6885), .O(n6897));
  orx   g06193(.a(n6872), .b(n6869), .O(n6898));
  andx  g06194(.a(n6864), .b(n6898), .O(n6899));
  orx   g06195(.a(n6873), .b(n6899), .O(n6900));
  orx   g06196(.a(n6886), .b(n6900), .O(n6901));
  orx   g06197(.a(n6882), .b(n6531), .O(n6902));
  orx   g06198(.a(n6878), .b(n6282), .O(n6903));
  andx  g06199(.a(n6903), .b(n6902), .O(n6904));
  orx   g06200(.a(n6886), .b(n6904), .O(n6905));
  andx  g06201(.a(n6905), .b(n6901), .O(n6906));
  andx  g06202(.a(n6906), .b(n6897), .O(n6907));
  andx  g06203(.a(n6907), .b(n6896), .O(n6908));
  invx  g06204(.a(n6908), .O(n6909));
  andx  g06205(.a(n6243), .b(n6211), .O(n6911));
  andx  g06206(.a(n6241), .b(n6224), .O(n6912));
  orx   g06207(.a(n6912), .b(n6911), .O(n6913));
  invx  g06208(.a(n6262), .O(n6914));
  andx  g06209(.a(n6619), .b(n6554), .O(n6916));
  orx   g06210(.a(n6916), .b(n6626), .O(n6917));
  orx   g06211(.a(n6917), .b(n6555), .O(n6918));
  orx   g06212(.a(n6262), .b(n6567), .O(n6920));
  andx  g06213(.a(n6920), .b(n6913), .O(n6921));
  andx  g06214(.a(n6914), .b(n6918), .O(n6924));
  andx  g06215(.a(n6924), .b(n6245), .O(n6925));
  orx   g06216(.a(n6925), .b(n6921), .O(n6926));
  andx  g06217(.a(n6926), .b(n6909), .O(n6927));
  orx   g06218(.a(n6924), .b(n6245), .O(n6929));
  orx   g06219(.a(n6920), .b(n6913), .O(n6930));
  andx  g06220(.a(n6930), .b(n6929), .O(n6931));
  andx  g06221(.a(n6931), .b(n6908), .O(n6932));
  orx   g06222(.a(n6932), .b(n6927), .O(n6933));
  orx   g06223(.a(n6608), .b(n6907), .O(n6936));
  andx  g06224(.a(n6936), .b(n6630), .O(n6937));
  andx  g06225(.a(n6609), .b(n6891), .O(n6940));
  andx  g06226(.a(n6940), .b(n6896), .O(n6941));
  orx   g06227(.a(n6941), .b(n6937), .O(n6942));
  andx  g06228(.a(n6886), .b(n6900), .O(n6951));
  orx   g06229(.a(n6951), .b(n6888), .O(n6952));
  orx   g06230(.a(n6952), .b(n6884), .O(n6953));
  orx   g06231(.a(n6887), .b(n6875), .O(n6954));
  andx  g06232(.a(n6954), .b(n6901), .O(n6955));
  orx   g06233(.a(n6955), .b(n6904), .O(n6956));
  andx  g06234(.a(n6956), .b(n6953), .O(n6957));
  andx  g06235(.a(n6655), .b(n6432), .O(n6961));
  andx  g06236(.a(n6651), .b(n6310), .O(n6962));
  orx   g06237(.a(n6962), .b(n6961), .O(n6963));
  invx  g06238(.a(n6807), .O(n6964));
  andx  g06239(.a(n6664), .b(n6329), .O(n6965));
  andx  g06240(.a(n6660), .b(n6435), .O(n6966));
  orx   g06241(.a(n6966), .b(n6965), .O(n6967));
  orx   g06242(.a(n6808), .b(n6967), .O(n6968));
  orx   g06243(.a(n6803), .b(n6792), .O(n6969));
  andx  g06244(.a(n6787), .b(n6969), .O(n6970));
  orx   g06245(.a(n6804), .b(n6970), .O(n6971));
  orx   g06246(.a(n6808), .b(n6971), .O(n6972));
  andx  g06247(.a(n6972), .b(n6968), .O(n6973));
  andx  g06248(.a(n6973), .b(n6964), .O(n6974));
  orx   g06249(.a(n6974), .b(n6963), .O(n6975));
  andx  g06250(.a(n6607), .b(n3645), .O(n6976));
  andx  g06251(.a(n6976), .b(n6975), .O(n6977));
  andx  g06252(.a(n6974), .b(n6963), .O(n6978));
  orx   g06253(.a(n6978), .b(n6977), .O(n6979));
  andx  g06254(.a(n6830), .b(n6979), .O(n6980));
  andx  g06255(.a(n6825), .b(n6819), .O(n6981));
  orx   g06256(.a(n6981), .b(n6980), .O(n6982));
  andx  g06257(.a(n6982), .b(n6824), .O(n6983));
  orx   g06258(.a(n6825), .b(n6819), .O(n6987));
  orx   g06259(.a(n6830), .b(n6979), .O(n6988));
  andx  g06260(.a(n6988), .b(n6987), .O(n6989));
  andx  g06261(.a(n6989), .b(n6648), .O(n6990));
  orx   g06262(.a(n6990), .b(n6983), .O(n6991));
  andx  g06263(.a(n165), .b(pi02), .O(n6992));
  andx  g06264(.a(n161), .b(pi03), .O(n6993));
  andx  g06265(.a(n103), .b(pi04), .O(n6994));
  andx  g06266(.a(pi19), .b(pi05), .O(n6995));
  orx   g06267(.a(n6995), .b(n6994), .O(n6996));
  orx   g06268(.a(n6996), .b(n6993), .O(n6997));
  orx   g06269(.a(n6997), .b(n6992), .O(n6998));
  andx  g06270(.a(n153), .b(pi01), .O(n6999));
  andx  g06271(.a(n148), .b(pi00), .O(n7000));
  orx   g06272(.a(n7000), .b(n6999), .O(n7001));
  orx   g06273(.a(n7001), .b(n6998), .O(n7002));
  andx  g06274(.a(n7002), .b(n3645), .O(n7003));
  invx  g06275(.a(n7003), .O(n7004));
  andx  g06276(.a(n7002), .b(n3180), .O(n7005));
  invx  g06277(.a(n7005), .O(n7006));
  orx   g06278(.a(n6730), .b(n6748), .O(n7007));
  orx   g06279(.a(n6740), .b(n6728), .O(n7008));
  andx  g06280(.a(n7008), .b(n7007), .O(n7009));
  orx   g06281(.a(n7009), .b(n6742), .O(n7010));
  andx  g06282(.a(n6740), .b(n6728), .O(n7011));
  andx  g06283(.a(n6730), .b(n6748), .O(n7012));
  orx   g06284(.a(n7012), .b(n7011), .O(n7013));
  orx   g06285(.a(n7013), .b(n6698), .O(n7014));
  andx  g06286(.a(n7014), .b(n7010), .O(n7015));
  andx  g06287(.a(n6726), .b(n6743), .O(n7016));
  orx   g06288(.a(n7016), .b(n6745), .O(n7017));
  invx  g06289(.a(n7017), .O(n7018));
  andx  g06290(.a(n7016), .b(n6745), .O(n7019));
  orx   g06291(.a(n7019), .b(n7018), .O(n7020));
  invx  g06292(.a(n6709), .O(n7021));
  andx  g06293(.a(n7021), .b(n6699), .O(n7022));
  invx  g06294(.a(n7022), .O(n7023));
  orx   g06295(.a(n7021), .b(n6699), .O(n7024));
  andx  g06296(.a(n7024), .b(n7023), .O(n7025));
  invx  g06297(.a(n6371), .O(n7026));
  orx   g06298(.a(n6370), .b(n6369), .O(n7027));
  andx  g06299(.a(n7027), .b(n7026), .O(n7028));
  andx  g06300(.a(n6704), .b(n7025), .O(n7030));
  invx  g06301(.a(n7030), .O(n7031));
  orx   g06302(.a(n6704), .b(n7025), .O(n7032));
  andx  g06303(.a(n7032), .b(n7031), .O(n7033));
  andx  g06304(.a(n7002), .b(n3258), .O(n7034));
  andx  g06305(.a(n7034), .b(n1790), .O(n7035));
  andx  g06306(.a(n7459), .b(n3230), .O(n7037));
  orx   g06307(.a(n6708), .b(n6707), .O(n7038));
  andx  g06308(.a(n7038), .b(n7021), .O(n7039));
  andx  g06309(.a(n7002), .b(n3230), .O(n7040));
  orx   g06310(.a(n7040), .b(n7459), .O(n7041));
  andx  g06311(.a(n7041), .b(n7039), .O(n7042));
  orx   g06312(.a(n7042), .b(n7037), .O(n7043));
  andx  g06313(.a(n7043), .b(n7033), .O(n7044));
  orx   g06314(.a(n7043), .b(n7033), .O(n7045));
  andx  g06315(.a(n7002), .b(n3221), .O(n7046));
  andx  g06316(.a(n7046), .b(n7045), .O(n7047));
  orx   g06317(.a(n7047), .b(n7044), .O(n7048));
  andx  g06318(.a(n7048), .b(n7020), .O(n7049));
  orx   g06319(.a(n7048), .b(n7020), .O(n7050));
  andx  g06320(.a(n7002), .b(n3210), .O(n7051));
  andx  g06321(.a(n7051), .b(n7050), .O(n7052));
  orx   g06322(.a(n7052), .b(n7049), .O(n7053));
  andx  g06323(.a(n7053), .b(n7015), .O(n7054));
  invx  g06324(.a(n7054), .O(n7055));
  andx  g06325(.a(n7013), .b(n6698), .O(n7056));
  andx  g06326(.a(n7009), .b(n6742), .O(n7057));
  orx   g06327(.a(n7057), .b(n7056), .O(n7058));
  invx  g06328(.a(n7049), .O(n7059));
  invx  g06329(.a(n7019), .O(n7060));
  andx  g06330(.a(n7060), .b(n7017), .O(n7061));
  invx  g06331(.a(n7048), .O(n7062));
  andx  g06332(.a(n7062), .b(n7061), .O(n7063));
  invx  g06333(.a(n7051), .O(n7064));
  orx   g06334(.a(n7064), .b(n7063), .O(n7065));
  andx  g06335(.a(n7065), .b(n7059), .O(n7066));
  andx  g06336(.a(n7066), .b(n7058), .O(n7067));
  andx  g06337(.a(n7002), .b(n3284), .O(n7068));
  invx  g06338(.a(n7068), .O(n7069));
  orx   g06339(.a(n7069), .b(n7067), .O(n7070));
  andx  g06340(.a(n7070), .b(n7055), .O(n7071));
  andx  g06341(.a(n7071), .b(n7006), .O(n7072));
  andx  g06342(.a(n6754), .b(n6733), .O(n7073));
  andx  g06343(.a(n6753), .b(n6751), .O(n7074));
  orx   g06344(.a(n7074), .b(n7073), .O(n7075));
  andx  g06345(.a(n7075), .b(n6738), .O(n7076));
  invx  g06346(.a(n7076), .O(n7077));
  orx   g06347(.a(n7075), .b(n6738), .O(n7078));
  andx  g06348(.a(n7078), .b(n7077), .O(n7079));
  orx   g06349(.a(n7079), .b(n7072), .O(n7080));
  orx   g06350(.a(n7071), .b(n3183), .O(n7081));
  andx  g06351(.a(n7081), .b(n7080), .O(n7082));
  andx  g06352(.a(n6759), .b(n6756), .O(n7083));
  andx  g06353(.a(n6758), .b(n6766), .O(n7084));
  orx   g06354(.a(n7084), .b(n7083), .O(n7085));
  andx  g06355(.a(n7085), .b(n6684), .O(n7086));
  orx   g06356(.a(n6758), .b(n6766), .O(n7087));
  orx   g06357(.a(n6759), .b(n6756), .O(n7088));
  andx  g06358(.a(n7088), .b(n7087), .O(n7089));
  andx  g06359(.a(n7089), .b(n6763), .O(n7090));
  orx   g06360(.a(n7090), .b(n7086), .O(n7091));
  andx  g06361(.a(n7091), .b(n7082), .O(n7092));
  andx  g06362(.a(n7002), .b(n3429), .O(n7093));
  invx  g06363(.a(n7093), .O(n7094));
  andx  g06364(.a(n7094), .b(n7082), .O(n7095));
  andx  g06365(.a(n7094), .b(n7091), .O(n7096));
  orx   g06366(.a(n7096), .b(n7095), .O(n7097));
  orx   g06367(.a(n7097), .b(n7092), .O(n7098));
  andx  g06368(.a(n7002), .b(n3171), .O(n7099));
  invx  g06369(.a(n7099), .O(n7100));
  andx  g06370(.a(n7100), .b(n7098), .O(n7101));
  andx  g06371(.a(n6781), .b(n6796), .O(n7105));
  andx  g06372(.a(n6780), .b(n6769), .O(n7106));
  orx   g06373(.a(n7106), .b(n7105), .O(n7107));
  andx  g06374(.a(n7107), .b(n6800), .O(n7108));
  orx   g06375(.a(n7107), .b(n6800), .O(n7109));
  invx  g06376(.a(n7109), .O(n7110));
  orx   g06377(.a(n7110), .b(n7108), .O(n7111));
  orx   g06378(.a(n7111), .b(n7101), .O(n7112));
  orx   g06379(.a(n7098), .b(n3418), .O(n7113));
  andx  g06380(.a(n7113), .b(n7112), .O(n7114));
  orx   g06381(.a(n6787), .b(n6785), .O(n7115));
  orx   g06382(.a(n6788), .b(n6803), .O(n7116));
  andx  g06383(.a(n7116), .b(n7115), .O(n7117));
  andx  g06384(.a(n7117), .b(n6675), .O(n7118));
  andx  g06385(.a(n6788), .b(n6803), .O(n7119));
  andx  g06386(.a(n6787), .b(n6785), .O(n7120));
  orx   g06387(.a(n7120), .b(n7119), .O(n7121));
  andx  g06388(.a(n7121), .b(n6792), .O(n7122));
  orx   g06389(.a(n7122), .b(n7118), .O(n7123));
  andx  g06390(.a(n7123), .b(n7114), .O(n7124));
  andx  g06391(.a(n7002), .b(n3413), .O(n7125));
  invx  g06392(.a(n7125), .O(n7126));
  andx  g06393(.a(n7126), .b(n7114), .O(n7127));
  andx  g06394(.a(n7126), .b(n7123), .O(n7128));
  orx   g06395(.a(n7128), .b(n7127), .O(n7129));
  orx   g06396(.a(n7129), .b(n7124), .O(n7130));
  andx  g06397(.a(n7130), .b(n7004), .O(n7131));
  andx  g06398(.a(n6808), .b(n6971), .O(n7132));
  orx   g06399(.a(n7132), .b(n6811), .O(n7133));
  orx   g06400(.a(n7133), .b(n6666), .O(n7134));
  invx  g06401(.a(n7134), .O(n7135));
  andx  g06402(.a(n7133), .b(n6666), .O(n7136));
  orx   g06403(.a(n7136), .b(n7135), .O(n7137));
  orx   g06404(.a(n7137), .b(n7131), .O(n7138));
  orx   g06405(.a(n7130), .b(n4509), .O(n7139));
  andx  g06406(.a(n7139), .b(n7138), .O(n7140));
  orx   g06407(.a(n6976), .b(n6813), .O(n7141));
  orx   g06408(.a(n6816), .b(n6974), .O(n7142));
  andx  g06409(.a(n7142), .b(n7141), .O(n7143));
  andx  g06410(.a(n7143), .b(n6657), .O(n7144));
  andx  g06411(.a(n6816), .b(n6974), .O(n7145));
  andx  g06412(.a(n6976), .b(n6813), .O(n7146));
  orx   g06413(.a(n7146), .b(n7145), .O(n7147));
  andx  g06414(.a(n7147), .b(n6963), .O(n7148));
  orx   g06415(.a(n7148), .b(n7144), .O(n7149));
  andx  g06416(.a(n7149), .b(n7140), .O(n7150));
  andx  g06417(.a(n7002), .b(n3721), .O(n7151));
  invx  g06418(.a(n7151), .O(n7152));
  andx  g06419(.a(n7152), .b(n7140), .O(n7153));
  andx  g06420(.a(n7152), .b(n7149), .O(n7154));
  orx   g06421(.a(n7154), .b(n7153), .O(n7155));
  orx   g06422(.a(n7155), .b(n7150), .O(n7156));
  orx   g06423(.a(n7156), .b(n6991), .O(n7157));
  andx  g06424(.a(n7002), .b(n4063), .O(n7158));
  invx  g06425(.a(n7158), .O(n7159));
  andx  g06426(.a(n7156), .b(n6991), .O(n7160));
  orx   g06427(.a(n7160), .b(n7159), .O(n7161));
  andx  g06428(.a(n7161), .b(n7157), .O(n7162));
  andx  g06429(.a(n6838), .b(n6844), .O(n7163));
  andx  g06430(.a(n6837), .b(n6834), .O(n7164));
  orx   g06431(.a(n7164), .b(n7163), .O(n7165));
  orx   g06432(.a(n7165), .b(n6639), .O(n7166));
  orx   g06433(.a(n6837), .b(n6834), .O(n7167));
  orx   g06434(.a(n6838), .b(n6844), .O(n7168));
  andx  g06435(.a(n7168), .b(n7167), .O(n7169));
  orx   g06436(.a(n7169), .b(n6841), .O(n7170));
  andx  g06437(.a(n7170), .b(n7166), .O(n7171));
  andx  g06438(.a(n7171), .b(n7162), .O(n7172));
  andx  g06439(.a(n7002), .b(n4114), .O(n7173));
  invx  g06440(.a(n7173), .O(n7174));
  orx   g06441(.a(n7174), .b(n7172), .O(n7175));
  orx   g06442(.a(n6989), .b(n6648), .O(n7176));
  orx   g06443(.a(n6982), .b(n6824), .O(n7177));
  andx  g06444(.a(n7177), .b(n7176), .O(n7178));
  invx  g06445(.a(n7150), .O(n7179));
  invx  g06446(.a(n7124), .O(n7180));
  invx  g06447(.a(n7092), .O(n7181));
  orx   g06448(.a(n7053), .b(n7015), .O(n7182));
  andx  g06449(.a(n7068), .b(n7182), .O(n7183));
  orx   g06450(.a(n7183), .b(n7054), .O(n7184));
  orx   g06451(.a(n7184), .b(n7005), .O(n7185));
  invx  g06452(.a(n7078), .O(n7186));
  orx   g06453(.a(n7186), .b(n7076), .O(n7187));
  andx  g06454(.a(n7187), .b(n7185), .O(n7188));
  andx  g06455(.a(n7184), .b(n3180), .O(n7189));
  orx   g06456(.a(n7189), .b(n7188), .O(n7190));
  orx   g06457(.a(n7093), .b(n7190), .O(n7191));
  orx   g06458(.a(n7089), .b(n6763), .O(n7192));
  orx   g06459(.a(n7085), .b(n6684), .O(n7193));
  andx  g06460(.a(n7193), .b(n7192), .O(n7194));
  orx   g06461(.a(n7093), .b(n7194), .O(n7195));
  andx  g06462(.a(n7195), .b(n7191), .O(n7196));
  andx  g06463(.a(n7196), .b(n7181), .O(n7197));
  orx   g06464(.a(n7099), .b(n7197), .O(n7198));
  invx  g06465(.a(n7108), .O(n7199));
  andx  g06466(.a(n7109), .b(n7199), .O(n7200));
  andx  g06467(.a(n7200), .b(n7198), .O(n7201));
  andx  g06468(.a(n7197), .b(n3171), .O(n7202));
  orx   g06469(.a(n7202), .b(n7201), .O(n7203));
  orx   g06470(.a(n7125), .b(n7203), .O(n7204));
  orx   g06471(.a(n7121), .b(n6792), .O(n7205));
  orx   g06472(.a(n7117), .b(n6675), .O(n7206));
  andx  g06473(.a(n7206), .b(n7205), .O(n7207));
  orx   g06474(.a(n7125), .b(n7207), .O(n7208));
  andx  g06475(.a(n7208), .b(n7204), .O(n7209));
  andx  g06476(.a(n7209), .b(n7180), .O(n7210));
  orx   g06477(.a(n7210), .b(n7003), .O(n7211));
  invx  g06478(.a(n7136), .O(n7212));
  andx  g06479(.a(n7212), .b(n7134), .O(n7213));
  andx  g06480(.a(n7213), .b(n7211), .O(n7214));
  andx  g06481(.a(n7210), .b(n3645), .O(n7215));
  orx   g06482(.a(n7215), .b(n7214), .O(n7216));
  orx   g06483(.a(n7151), .b(n7216), .O(n7217));
  orx   g06484(.a(n7147), .b(n6963), .O(n7218));
  orx   g06485(.a(n7143), .b(n6657), .O(n7219));
  andx  g06486(.a(n7219), .b(n7218), .O(n7220));
  orx   g06487(.a(n7151), .b(n7220), .O(n7221));
  andx  g06488(.a(n7221), .b(n7217), .O(n7222));
  andx  g06489(.a(n7222), .b(n7179), .O(n7223));
  andx  g06490(.a(n7223), .b(n7178), .O(n7224));
  orx   g06491(.a(n7223), .b(n7178), .O(n7225));
  andx  g06492(.a(n7225), .b(n7158), .O(n7226));
  orx   g06493(.a(n7226), .b(n7224), .O(n7227));
  andx  g06494(.a(n7169), .b(n6841), .O(n7228));
  andx  g06495(.a(n7165), .b(n6639), .O(n7229));
  orx   g06496(.a(n7229), .b(n7228), .O(n7230));
  andx  g06497(.a(n7230), .b(n7227), .O(n7231));
  invx  g06498(.a(n7231), .O(n7232));
  andx  g06499(.a(n7232), .b(n7175), .O(n7233));
  orx   g06500(.a(n6864), .b(n6847), .O(n7234));
  orx   g06501(.a(n6865), .b(n6869), .O(n7235));
  andx  g06502(.a(n7235), .b(n7234), .O(n7236));
  andx  g06503(.a(n7236), .b(n6862), .O(n7237));
  andx  g06504(.a(n6865), .b(n6869), .O(n7238));
  andx  g06505(.a(n6864), .b(n6847), .O(n7239));
  orx   g06506(.a(n7239), .b(n7238), .O(n7240));
  andx  g06507(.a(n7240), .b(n6872), .O(n7241));
  orx   g06508(.a(n7241), .b(n7237), .O(n7242));
  andx  g06509(.a(n7242), .b(n7233), .O(n7243));
  invx  g06510(.a(n7243), .O(n7244));
  orx   g06511(.a(n7230), .b(n7227), .O(n7245));
  andx  g06512(.a(n7173), .b(n7245), .O(n7246));
  orx   g06513(.a(n7231), .b(n7246), .O(n7247));
  andx  g06514(.a(n7002), .b(n4490), .O(n7248));
  orx   g06515(.a(n7248), .b(n7247), .O(n7249));
  orx   g06516(.a(n7240), .b(n6872), .O(n7250));
  orx   g06517(.a(n7236), .b(n6862), .O(n7251));
  andx  g06518(.a(n7251), .b(n7250), .O(n7252));
  orx   g06519(.a(n7248), .b(n7252), .O(n7253));
  andx  g06520(.a(n7253), .b(n7249), .O(n7254));
  andx  g06521(.a(n7254), .b(n7244), .O(n7255));
  andx  g06522(.a(n7002), .b(n2724), .O(n7257));
  andx  g06523(.a(n7255), .b(n6957), .O(n7259));
  andx  g06524(.a(n7259), .b(n6942), .O(n7261));
  invx  g06525(.a(n6568), .O(n7262));
  andx  g06526(.a(n7262), .b(n6240), .O(n7263));
  andx  g06527(.a(n6237), .b(n6234), .O(n7264));
  orx   g06528(.a(n6573), .b(n7264), .O(n7266));
  andx  g06529(.a(n6568), .b(n7266), .O(n7267));
  orx   g06530(.a(n7267), .b(n7263), .O(n7268));
  andx  g06531(.a(n6926), .b(n6908), .O(n7269));
  orx   g06532(.a(n7269), .b(n7268), .O(n7270));
  andx  g06533(.a(n7269), .b(n7268), .O(n7273));
  andx  g06534(.a(n6593), .b(n6572), .O(n7276));
  andx  g06535(.a(n6587), .b(n6573), .O(n7277));
  orx   g06536(.a(n7277), .b(n7276), .O(n7278));
  invx  g06537(.a(n5771), .O(n7280));
  andx  g06538(.a(n7280), .b(n5407), .O(n7281));
  orx   g06539(.a(n5368), .b(n5403), .O(n7282));
  orx   g06540(.a(n5398), .b(n5378), .O(n7283));
  andx  g06541(.a(n7283), .b(n7282), .O(n7284));
  andx  g06542(.a(n5771), .b(n7284), .O(n7285));
  orx   g06543(.a(n7285), .b(n7281), .O(n7286));
  orx   g06544(.a(n6940), .b(n6896), .O(n7288));
  orx   g06545(.a(n6936), .b(n6630), .O(n7289));
  andx  g06546(.a(n7289), .b(n7288), .O(n7290));
  andx  g06547(.a(n6955), .b(n6904), .O(n7291));
  andx  g06548(.a(n6952), .b(n6884), .O(n7292));
  orx   g06549(.a(n7292), .b(n7291), .O(n7293));
  invx  g06550(.a(n7248), .O(n7294));
  andx  g06551(.a(n7294), .b(n7233), .O(n7295));
  andx  g06552(.a(n7294), .b(n7242), .O(n7296));
  orx   g06553(.a(n7296), .b(n7295), .O(n7297));
  orx   g06554(.a(n7297), .b(n7243), .O(n7298));
  invx  g06555(.a(n7257), .O(n7300));
  andx  g06556(.a(n7310), .b(n7290), .O(n7304));
  invx  g06557(.a(n7304), .O(n7305));
  orx   g06558(.a(n7310), .b(n7290), .O(n7306));
  andx  g06559(.a(n7300), .b(n7298), .O(n7308));
  orx   g06560(.a(n7308), .b(n7293), .O(n7310));
  orx   g06561(.a(n7257), .b(n7255), .O(n7312));
  orx   g06562(.a(n7312), .b(n6957), .O(n7314));
  andx  g06563(.a(n7314), .b(n7310), .O(n7315));
  orx   g06564(.a(n7294), .b(n7233), .O(n7323));
  andx  g06565(.a(n7323), .b(n7249), .O(n7324));
  andx  g06566(.a(n7324), .b(n7252), .O(n7325));
  andx  g06567(.a(n7248), .b(n7247), .O(n7328));
  orx   g06568(.a(n7328), .b(n7295), .O(n7329));
  andx  g06569(.a(n7329), .b(n7242), .O(n7330));
  orx   g06570(.a(n7330), .b(n7325), .O(n7331));
  orx   g06571(.a(n7173), .b(n7162), .O(n7332));
  orx   g06572(.a(n7174), .b(n7227), .O(n7333));
  andx  g06573(.a(n7333), .b(n7332), .O(n7334));
  orx   g06574(.a(n7334), .b(n7230), .O(n7335));
  andx  g06575(.a(n7174), .b(n7227), .O(n7336));
  andx  g06576(.a(n7173), .b(n7162), .O(n7337));
  orx   g06577(.a(n7337), .b(n7336), .O(n7338));
  orx   g06578(.a(n7338), .b(n7171), .O(n7339));
  andx  g06579(.a(n7339), .b(n7335), .O(n7340));
  andx  g06580(.a(n7151), .b(n7216), .O(n7349));
  orx   g06581(.a(n7349), .b(n7153), .O(n7350));
  andx  g06582(.a(n7350), .b(n7220), .O(n7351));
  orx   g06583(.a(n7152), .b(n7140), .O(n7352));
  andx  g06584(.a(n7352), .b(n7217), .O(n7353));
  andx  g06585(.a(n7353), .b(n7149), .O(n7354));
  orx   g06586(.a(n7354), .b(n7351), .O(n7355));
  andx  g06587(.a(n153), .b(pi00), .O(n7356));
  andx  g06588(.a(n165), .b(pi01), .O(n7357));
  andx  g06589(.a(n161), .b(pi02), .O(n7358));
  andx  g06590(.a(n103), .b(pi03), .O(n7359));
  andx  g06591(.a(pi19), .b(pi04), .O(n7360));
  orx   g06592(.a(n7360), .b(n7359), .O(n7361));
  orx   g06593(.a(n7361), .b(n7358), .O(n7362));
  orx   g06594(.a(n7362), .b(n7357), .O(n7363));
  orx   g06595(.a(n7363), .b(n7356), .O(n7364));
  andx  g06596(.a(n7364), .b(n3721), .O(n7365));
  andx  g06597(.a(n7139), .b(n7211), .O(n7366));
  orx   g06598(.a(n7366), .b(n7213), .O(n7367));
  orx   g06599(.a(n7215), .b(n7131), .O(n7368));
  orx   g06600(.a(n7368), .b(n7137), .O(n7369));
  andx  g06601(.a(n7369), .b(n7367), .O(n7370));
  andx  g06602(.a(n7370), .b(n7365), .O(n7371));
  andx  g06603(.a(n7364), .b(n3645), .O(n7372));
  andx  g06604(.a(n7125), .b(n7203), .O(n7381));
  orx   g06605(.a(n7381), .b(n7127), .O(n7382));
  andx  g06606(.a(n7382), .b(n7207), .O(n7383));
  orx   g06607(.a(n7126), .b(n7114), .O(n7384));
  andx  g06608(.a(n7384), .b(n7204), .O(n7385));
  andx  g06609(.a(n7385), .b(n7123), .O(n7386));
  orx   g06610(.a(n7386), .b(n7383), .O(n7387));
  andx  g06611(.a(n7387), .b(n7372), .O(n7388));
  andx  g06612(.a(n7364), .b(n3171), .O(n7389));
  andx  g06613(.a(n7093), .b(n7190), .O(n7397));
  orx   g06614(.a(n7397), .b(n7095), .O(n7398));
  andx  g06615(.a(n7398), .b(n7194), .O(n7399));
  orx   g06616(.a(n7094), .b(n7082), .O(n7401));
  andx  g06617(.a(n7401), .b(n7191), .O(n7402));
  andx  g06618(.a(n7402), .b(n7091), .O(n7403));
  orx   g06619(.a(n7403), .b(n7399), .O(n7404));
  andx  g06620(.a(n7404), .b(n7389), .O(n7405));
  orx   g06621(.a(n7069), .b(n7066), .O(n7406));
  orx   g06622(.a(n7068), .b(n7053), .O(n7407));
  andx  g06623(.a(n7407), .b(n7406), .O(n7408));
  orx   g06624(.a(n7408), .b(n7015), .O(n7409));
  andx  g06625(.a(n7068), .b(n7053), .O(n7410));
  andx  g06626(.a(n7069), .b(n7066), .O(n7411));
  orx   g06627(.a(n7411), .b(n7410), .O(n7412));
  orx   g06628(.a(n7412), .b(n7058), .O(n7413));
  andx  g06629(.a(n7413), .b(n7409), .O(n7414));
  andx  g06630(.a(n7364), .b(n3180), .O(n7415));
  andx  g06631(.a(n7415), .b(n7414), .O(n7416));
  andx  g06632(.a(n7064), .b(n7048), .O(n7417));
  invx  g06633(.a(n7417), .O(n7418));
  orx   g06634(.a(n7064), .b(n7048), .O(n7419));
  andx  g06635(.a(n7419), .b(n7418), .O(n7420));
  orx   g06636(.a(n7420), .b(n7061), .O(n7421));
  invx  g06637(.a(n7419), .O(n7422));
  orx   g06638(.a(n7422), .b(n7417), .O(n7423));
  orx   g06639(.a(n7423), .b(n7020), .O(n7424));
  andx  g06640(.a(n7424), .b(n7421), .O(n7425));
  invx  g06641(.a(n7043), .O(n7426));
  andx  g06642(.a(n7046), .b(n7426), .O(n7427));
  invx  g06643(.a(n7427), .O(n7428));
  orx   g06644(.a(n7046), .b(n7426), .O(n7429));
  andx  g06645(.a(n7429), .b(n7428), .O(n7430));
  invx  g06646(.a(n7430), .O(n7431));
  andx  g06647(.a(n7431), .b(n7033), .O(n7432));
  orx   g06648(.a(n7431), .b(n7033), .O(n7433));
  invx  g06649(.a(n7433), .O(n7434));
  orx   g06650(.a(n7434), .b(n7432), .O(n7435));
  andx  g06651(.a(n7364), .b(n3210), .O(n7436));
  invx  g06652(.a(n7436), .O(n7437));
  andx  g06653(.a(n7437), .b(n7435), .O(n7438));
  invx  g06654(.a(n7438), .O(n7439));
  invx  g06655(.a(n7432), .O(n7440));
  andx  g06656(.a(n7433), .b(n7440), .O(n7441));
  andx  g06657(.a(n7436), .b(n7441), .O(n7442));
  invx  g06658(.a(n7039), .O(n7443));
  invx  g06659(.a(n7037), .O(n7444));
  andx  g06660(.a(n7041), .b(n7444), .O(n7445));
  invx  g06661(.a(n7445), .O(n7446));
  andx  g06662(.a(n7446), .b(n7443), .O(n7447));
  andx  g06663(.a(n7445), .b(n7039), .O(n7448));
  orx   g06664(.a(n7448), .b(n7447), .O(n7449));
  invx  g06665(.a(n7449), .O(n7450));
  andx  g06666(.a(n7364), .b(n3221), .O(n7451));
  andx  g06667(.a(n7451), .b(n7450), .O(n7452));
  invx  g06668(.a(n7452), .O(n7453));
  andx  g06669(.a(n7449), .b(n3236), .O(n7454));
  invx  g06670(.a(n7034), .O(n7455));
  andx  g06671(.a(n6607), .b(n1790), .O(n7456));
  invx  g06672(.a(n7456), .O(n7457));
  andx  g06673(.a(n7457), .b(n7455), .O(n7458));
  andx  g06674(.a(n7456), .b(n7034), .O(n7459));
  orx   g06675(.a(n7459), .b(n7458), .O(n7460));
  invx  g06676(.a(n7460), .O(n7461));
  andx  g06677(.a(n7461), .b(n7035), .O(n7462));
  orx   g06678(.a(n7462), .b(n3230), .O(n7463));
  orx   g06679(.a(n7461), .b(n7035), .O(n7464));
  andx  g06680(.a(n7464), .b(n7364), .O(n7465));
  andx  g06681(.a(n7465), .b(n7463), .O(n7466));
  invx  g06682(.a(n7466), .O(n7467));
  orx   g06683(.a(n7467), .b(n7454), .O(n7468));
  andx  g06684(.a(n7468), .b(n7453), .O(n7469));
  invx  g06685(.a(n7469), .O(n7470));
  orx   g06686(.a(n7470), .b(n7442), .O(n7471));
  andx  g06687(.a(n7471), .b(n7439), .O(n7472));
  andx  g06688(.a(n7472), .b(n7425), .O(n7473));
  orx   g06689(.a(n7472), .b(n7425), .O(n7474));
  andx  g06690(.a(n7364), .b(n3284), .O(n7475));
  andx  g06691(.a(n7475), .b(n7474), .O(n7476));
  orx   g06692(.a(n7476), .b(n7473), .O(n7477));
  andx  g06693(.a(n7477), .b(n7414), .O(n7478));
  andx  g06694(.a(n7477), .b(n7415), .O(n7479));
  orx   g06695(.a(n7479), .b(n7478), .O(n7480));
  orx   g06696(.a(n7480), .b(n7416), .O(n7481));
  orx   g06697(.a(n7189), .b(n7072), .O(n7482));
  andx  g06698(.a(n7482), .b(n7187), .O(n7483));
  andx  g06699(.a(n7081), .b(n7185), .O(n7484));
  andx  g06700(.a(n7484), .b(n7079), .O(n7485));
  orx   g06701(.a(n7485), .b(n7483), .O(n7486));
  andx  g06702(.a(n7486), .b(n7481), .O(n7487));
  orx   g06703(.a(n7486), .b(n7481), .O(n7491));
  andx  g06704(.a(n7364), .b(n3429), .O(n7492));
  andx  g06705(.a(n7492), .b(n7491), .O(n7493));
  orx   g06706(.a(n7493), .b(n7487), .O(n7494));
  andx  g06707(.a(n7494), .b(n7389), .O(n7495));
  andx  g06708(.a(n7494), .b(n7404), .O(n7496));
  orx   g06709(.a(n7496), .b(n7495), .O(n7497));
  orx   g06710(.a(n7497), .b(n7405), .O(n7498));
  orx   g06711(.a(n7202), .b(n7101), .O(n7499));
  andx  g06712(.a(n7499), .b(n7200), .O(n7500));
  andx  g06713(.a(n7113), .b(n7198), .O(n7501));
  andx  g06714(.a(n7501), .b(n7111), .O(n7502));
  orx   g06715(.a(n7502), .b(n7500), .O(n7503));
  andx  g06716(.a(n7503), .b(n7498), .O(n7504));
  orx   g06717(.a(n7503), .b(n7498), .O(n7508));
  andx  g06718(.a(n7364), .b(n3413), .O(n7509));
  andx  g06719(.a(n7509), .b(n7508), .O(n7510));
  orx   g06720(.a(n7510), .b(n7504), .O(n7511));
  andx  g06721(.a(n7511), .b(n7372), .O(n7512));
  andx  g06722(.a(n7511), .b(n7387), .O(n7513));
  orx   g06723(.a(n7513), .b(n7512), .O(n7514));
  orx   g06724(.a(n7514), .b(n7388), .O(n7515));
  andx  g06725(.a(n7515), .b(n7365), .O(n7516));
  andx  g06726(.a(n7515), .b(n7370), .O(n7517));
  orx   g06727(.a(n7517), .b(n7516), .O(n7518));
  orx   g06728(.a(n7518), .b(n7371), .O(n7519));
  andx  g06729(.a(n7519), .b(n7355), .O(n7520));
  andx  g06730(.a(n7364), .b(n4063), .O(n7521));
  andx  g06731(.a(n7521), .b(n7355), .O(n7522));
  andx  g06732(.a(n7521), .b(n7519), .O(n7523));
  orx   g06733(.a(n7523), .b(n7522), .O(n7524));
  orx   g06734(.a(n7524), .b(n7520), .O(n7525));
  orx   g06735(.a(n7158), .b(n7223), .O(n7526));
  orx   g06736(.a(n7159), .b(n7156), .O(n7527));
  andx  g06737(.a(n7527), .b(n7526), .O(n7528));
  andx  g06738(.a(n7528), .b(n6991), .O(n7529));
  andx  g06739(.a(n7159), .b(n7156), .O(n7530));
  andx  g06740(.a(n7158), .b(n7223), .O(n7531));
  orx   g06741(.a(n7531), .b(n7530), .O(n7532));
  andx  g06742(.a(n7532), .b(n7178), .O(n7533));
  orx   g06743(.a(n7533), .b(n7529), .O(n7534));
  andx  g06744(.a(n7534), .b(n7525), .O(n7535));
  invx  g06745(.a(n7535), .O(n7536));
  invx  g06746(.a(n7520), .O(n7537));
  orx   g06747(.a(n7353), .b(n7149), .O(n7538));
  orx   g06748(.a(n7350), .b(n7220), .O(n7539));
  andx  g06749(.a(n7539), .b(n7538), .O(n7540));
  invx  g06750(.a(n7521), .O(n7541));
  orx   g06751(.a(n7541), .b(n7540), .O(n7542));
  invx  g06752(.a(n7371), .O(n7543));
  invx  g06753(.a(n7365), .O(n7544));
  invx  g06754(.a(n7388), .O(n7545));
  invx  g06755(.a(n7372), .O(n7546));
  invx  g06756(.a(n7504), .O(n7547));
  invx  g06757(.a(n7405), .O(n7548));
  invx  g06758(.a(n7389), .O(n7549));
  invx  g06759(.a(n7487), .O(n7550));
  invx  g06760(.a(n7416), .O(n7551));
  andx  g06761(.a(n7412), .b(n7058), .O(n7552));
  andx  g06762(.a(n7408), .b(n7015), .O(n7553));
  orx   g06763(.a(n7553), .b(n7552), .O(n7554));
  invx  g06764(.a(n7473), .O(n7555));
  andx  g06765(.a(n7423), .b(n7020), .O(n7556));
  andx  g06766(.a(n7420), .b(n7061), .O(n7557));
  orx   g06767(.a(n7557), .b(n7556), .O(n7558));
  orx   g06768(.a(n7437), .b(n7435), .O(n7559));
  andx  g06769(.a(n7469), .b(n7559), .O(n7560));
  orx   g06770(.a(n7560), .b(n7438), .O(n7561));
  andx  g06771(.a(n7561), .b(n7558), .O(n7562));
  invx  g06772(.a(n7475), .O(n7563));
  orx   g06773(.a(n7563), .b(n7562), .O(n7564));
  andx  g06774(.a(n7564), .b(n7555), .O(n7565));
  orx   g06775(.a(n7565), .b(n7554), .O(n7566));
  invx  g06776(.a(n7415), .O(n7567));
  orx   g06777(.a(n7565), .b(n7567), .O(n7568));
  andx  g06778(.a(n7568), .b(n7566), .O(n7569));
  andx  g06779(.a(n7569), .b(n7551), .O(n7570));
  andx  g06780(.a(n7482), .b(n7079), .O(n7571));
  andx  g06781(.a(n7484), .b(n7187), .O(n7572));
  orx   g06782(.a(n7572), .b(n7571), .O(n7573));
  andx  g06783(.a(n7573), .b(n7570), .O(n7574));
  invx  g06784(.a(n7492), .O(n7575));
  orx   g06785(.a(n7575), .b(n7574), .O(n7576));
  andx  g06786(.a(n7576), .b(n7550), .O(n7577));
  orx   g06787(.a(n7577), .b(n7549), .O(n7578));
  orx   g06788(.a(n7402), .b(n7091), .O(n7579));
  orx   g06789(.a(n7398), .b(n7194), .O(n7580));
  andx  g06790(.a(n7580), .b(n7579), .O(n7581));
  orx   g06791(.a(n7577), .b(n7581), .O(n7582));
  andx  g06792(.a(n7582), .b(n7578), .O(n7583));
  andx  g06793(.a(n7583), .b(n7548), .O(n7584));
  andx  g06794(.a(n7499), .b(n7111), .O(n7585));
  andx  g06795(.a(n7501), .b(n7200), .O(n7586));
  orx   g06796(.a(n7586), .b(n7585), .O(n7587));
  andx  g06797(.a(n7587), .b(n7584), .O(n7588));
  invx  g06798(.a(n7509), .O(n7589));
  orx   g06799(.a(n7589), .b(n7588), .O(n7590));
  andx  g06800(.a(n7590), .b(n7547), .O(n7591));
  orx   g06801(.a(n7591), .b(n7546), .O(n7592));
  orx   g06802(.a(n7385), .b(n7123), .O(n7593));
  orx   g06803(.a(n7382), .b(n7207), .O(n7594));
  andx  g06804(.a(n7594), .b(n7593), .O(n7595));
  orx   g06805(.a(n7591), .b(n7595), .O(n7596));
  andx  g06806(.a(n7596), .b(n7592), .O(n7597));
  andx  g06807(.a(n7597), .b(n7545), .O(n7598));
  orx   g06808(.a(n7598), .b(n7544), .O(n7599));
  andx  g06809(.a(n7368), .b(n7137), .O(n7600));
  andx  g06810(.a(n7366), .b(n7213), .O(n7601));
  orx   g06811(.a(n7601), .b(n7600), .O(n7602));
  orx   g06812(.a(n7598), .b(n7602), .O(n7603));
  andx  g06813(.a(n7603), .b(n7599), .O(n7604));
  andx  g06814(.a(n7604), .b(n7543), .O(n7605));
  orx   g06815(.a(n7541), .b(n7605), .O(n7606));
  andx  g06816(.a(n7606), .b(n7542), .O(n7607));
  andx  g06817(.a(n7607), .b(n7537), .O(n7608));
  orx   g06818(.a(n7532), .b(n7178), .O(n7609));
  orx   g06819(.a(n7528), .b(n6991), .O(n7610));
  andx  g06820(.a(n7610), .b(n7609), .O(n7611));
  andx  g06821(.a(n7611), .b(n7608), .O(n7612));
  andx  g06822(.a(n7364), .b(n4114), .O(n7613));
  invx  g06823(.a(n7613), .O(n7614));
  orx   g06824(.a(n7614), .b(n7612), .O(n7615));
  andx  g06825(.a(n7615), .b(n7536), .O(n7616));
  andx  g06826(.a(n7616), .b(n7340), .O(n7617));
  andx  g06827(.a(n7364), .b(n4490), .O(n7618));
  invx  g06828(.a(n7618), .O(n7619));
  orx   g06829(.a(n7619), .b(n7617), .O(n7620));
  orx   g06830(.a(n7616), .b(n7340), .O(n7621));
  andx  g06831(.a(n7621), .b(n7620), .O(n7622));
  andx  g06832(.a(n7364), .b(n2724), .O(n7624));
  invx  g06833(.a(n7624), .O(n7625));
  orx   g06834(.a(n7329), .b(n7242), .O(n7627));
  orx   g06835(.a(n7324), .b(n7252), .O(n7628));
  andx  g06836(.a(n7628), .b(n7627), .O(n7629));
  andx  g06837(.a(n7338), .b(n7171), .O(n7630));
  andx  g06838(.a(n7334), .b(n7230), .O(n7631));
  orx   g06839(.a(n7631), .b(n7630), .O(n7632));
  orx   g06840(.a(n7534), .b(n7525), .O(n7633));
  andx  g06841(.a(n7613), .b(n7633), .O(n7634));
  orx   g06842(.a(n7634), .b(n7535), .O(n7635));
  orx   g06843(.a(n7635), .b(n7632), .O(n7636));
  andx  g06844(.a(n7618), .b(n7636), .O(n7637));
  andx  g06845(.a(n7635), .b(n7632), .O(n7638));
  orx   g06846(.a(n7638), .b(n7637), .O(n7639));
  andx  g06847(.a(n7639), .b(n7629), .O(n7640));
  invx  g06848(.a(n7640), .O(n7641));
  andx  g06849(.a(n7640), .b(n7315), .O(n7644));
  andx  g06850(.a(n7644), .b(n7305), .O(n7646));
  andx  g06851(.a(n5866), .b(n5397), .O(n7652));
  andx  g06852(.a(n7652), .b(n5781), .O(n7653));
  andx  g06853(.a(n7653), .b(n5390), .O(n7654));
  andx  g06854(.a(n7654), .b(n7868), .O(n7655));
  orx   g06855(.a(n7655), .b(n5867), .O(n7656));
  invx  g06856(.a(n7656), .O(n7657));
  andx  g06857(.a(n5858), .b(n5863), .O(n7658));
  invx  g06858(.a(n7658), .O(n7659));
  andx  g06859(.a(n5845), .b(n5853), .O(n7660));
  orx   g06860(.a(n7660), .b(n5846), .O(n7661));
  invx  g06861(.a(n7661), .O(n7662));
  andx  g06862(.a(n4114), .b(n299), .O(n7663));
  andx  g06863(.a(n5811), .b(n5792), .O(n7664));
  invx  g06864(.a(n7664), .O(n7665));
  andx  g06865(.a(n5810), .b(n5789), .O(n7666));
  orx   g06866(.a(n7666), .b(n5793), .O(n7667));
  andx  g06867(.a(n7667), .b(n7665), .O(n7668));
  invx  g06868(.a(n7668), .O(n7669));
  andx  g06869(.a(n7669), .b(n7663), .O(n7670));
  invx  g06870(.a(n7663), .O(n7671));
  andx  g06871(.a(n7668), .b(n7671), .O(n7672));
  orx   g06872(.a(n7672), .b(n7670), .O(n7673));
  invx  g06873(.a(n7673), .O(n7674));
  andx  g06874(.a(n4063), .b(n827), .O(n7675));
  invx  g06875(.a(n7675), .O(n7676));
  andx  g06876(.a(n7676), .b(n3721), .O(n7677));
  andx  g06877(.a(n6829), .b(n827), .O(n7678));
  andx  g06878(.a(n7678), .b(n4063), .O(n7679));
  orx   g06879(.a(n7679), .b(n7677), .O(n7680));
  andx  g06880(.a(n5806), .b(n5799), .O(n7681));
  orx   g06881(.a(n7681), .b(n4509), .O(n7682));
  orx   g06882(.a(n5806), .b(n6829), .O(n7683));
  andx  g06883(.a(n7683), .b(n7682), .O(n7684));
  invx  g06884(.a(n7684), .O(n7685));
  andx  g06885(.a(n7685), .b(n7680), .O(n7686));
  invx  g06886(.a(n7686), .O(n7687));
  orx   g06887(.a(n7685), .b(n7680), .O(n7688));
  andx  g06888(.a(n7688), .b(n7687), .O(n7689));
  andx  g06889(.a(n7689), .b(n7674), .O(n7690));
  invx  g06890(.a(n7689), .O(n7691));
  andx  g06891(.a(n7691), .b(n7673), .O(n7692));
  orx   g06892(.a(n7692), .b(n7690), .O(n7693));
  andx  g06893(.a(n5822), .b(n5815), .O(n7694));
  orx   g06894(.a(n7694), .b(n5819), .O(n7695));
  invx  g06895(.a(n7695), .O(n7697));
  andx  g06896(.a(n338), .b(n7697), .O(n7700));
  invx  g06897(.a(n7700), .O(n7701));
  andx  g06898(.a(n7701), .b(n7693), .O(n7702));
  invx  g06899(.a(n7693), .O(n7703));
  andx  g06900(.a(n7700), .b(n7703), .O(n7704));
  orx   g06901(.a(n7704), .b(n7702), .O(n7705));
  invx  g06902(.a(n7705), .O(n7706));
  andx  g06903(.a(n2724), .b(n376), .O(n7707));
  andx  g06904(.a(n5835), .b(n5827), .O(n7708));
  orx   g06905(.a(n7708), .b(n467), .O(n7709));
  invx  g06906(.a(n7709), .O(n7712));
  andx  g06907(.a(n7712), .b(n7706), .O(n7718));
  andx  g06908(.a(n7709), .b(n7705), .O(n7719));
  orx   g06909(.a(n7719), .b(n7718), .O(n7720));
  invx  g06910(.a(n7720), .O(n7721));
  andx  g06911(.a(n7721), .b(n7662), .O(n7722));
  andx  g06912(.a(n7720), .b(n7661), .O(n7723));
  orx   g06913(.a(n7723), .b(n7722), .O(n7724));
  andx  g06914(.a(n7724), .b(n7659), .O(n7725));
  andx  g06915(.a(n7725), .b(n7657), .O(n7726));
  invx  g06916(.a(n7724), .O(n7727));
  andx  g06917(.a(n7727), .b(n7658), .O(n7728));
  andx  g06918(.a(n7727), .b(n7656), .O(n7729));
  orx   g06919(.a(n7729), .b(n7728), .O(n7730));
  orx   g06920(.a(n7730), .b(n7726), .O(n7731));
  invx  g06921(.a(n7731), .O(n7732));
  invx  g06922(.a(n5390), .O(n7733));
  orx   g06923(.a(n7733), .b(n5389), .O(n7734));
  orx   g06924(.a(n5395), .b(n5088), .O(n7735));
  orx   g06925(.a(n5381), .b(n5393), .O(n7736));
  andx  g06926(.a(n7736), .b(n7735), .O(n7737));
  invx  g06927(.a(n5777), .O(n7738));
  invx  g06928(.a(n7644), .O(n7740));
  orx   g06929(.a(n7740), .b(n7304), .O(n7742));
  orx   g06930(.a(n6568), .b(n7266), .O(n7743));
  orx   g06931(.a(n7262), .b(n6240), .O(n7744));
  andx  g06932(.a(n7744), .b(n7743), .O(n7745));
  invx  g06933(.a(n7269), .O(n7746));
  andx  g06934(.a(n7746), .b(n7745), .O(n7747));
  andx  g06935(.a(n7869), .b(n7738), .O(n7756));
  orx   g06936(.a(n7756), .b(n7737), .O(n7757));
  andx  g06937(.a(n7757), .b(n7734), .O(n7758));
  invx  g06938(.a(n5389), .O(n7759));
  andx  g06939(.a(n5390), .b(n7759), .O(n7760));
  invx  g06940(.a(n7757), .O(n7761));
  orx   g06941(.a(n7882), .b(n7758), .O(n7763));
  orx   g06942(.a(n7746), .b(n7745), .O(n7764));
  andx  g06943(.a(n7764), .b(n7270), .O(n7765));
  orx   g06944(.a(n6931), .b(n6908), .O(n7766));
  orx   g06945(.a(n6926), .b(n6909), .O(n7767));
  andx  g06946(.a(n7767), .b(n7766), .O(n7768));
  andx  g06947(.a(n7742), .b(n7306), .O(n7769));
  orx   g06948(.a(n7769), .b(n7768), .O(n7770));
  orx   g06949(.a(n7770), .b(n7765), .O(n7771));
  orx   g06950(.a(n7273), .b(n7747), .O(n7772));
  invx  g06951(.a(n7770), .O(n7773));
  orx   g06952(.a(n7773), .b(n7772), .O(n7774));
  andx  g06953(.a(n7774), .b(n7771), .O(n7775));
  andx  g06954(.a(n7613), .b(n7608), .O(n7776));
  andx  g06955(.a(n7614), .b(n7525), .O(n7777));
  orx   g06956(.a(n7777), .b(n7776), .O(n7778));
  orx   g06957(.a(n7778), .b(n7611), .O(n7779));
  orx   g06958(.a(n7614), .b(n7525), .O(n7780));
  orx   g06959(.a(n7613), .b(n7608), .O(n7781));
  andx  g06960(.a(n7781), .b(n7780), .O(n7782));
  orx   g06961(.a(n7782), .b(n7534), .O(n7783));
  andx  g06962(.a(n7783), .b(n7779), .O(n7784));
  andx  g06963(.a(n7515), .b(n7544), .O(n7785));
  andx  g06964(.a(n7598), .b(n7365), .O(n7786));
  orx   g06965(.a(n7786), .b(n7785), .O(n7787));
  invx  g06966(.a(n7787), .O(n7788));
  andx  g06967(.a(n7788), .b(n7370), .O(n7789));
  andx  g06968(.a(n7787), .b(n7602), .O(n7790));
  orx   g06969(.a(n7790), .b(n7789), .O(n7791));
  invx  g06970(.a(n7791), .O(n7792));
  andx  g06971(.a(n7521), .b(n7605), .O(n7800));
  andx  g06972(.a(n7541), .b(n7519), .O(n7801));
  orx   g06973(.a(n7801), .b(n7800), .O(n7802));
  orx   g06974(.a(n7802), .b(n7355), .O(n7803));
  invx  g06975(.a(n7803), .O(n7804));
  andx  g06976(.a(n7802), .b(n7355), .O(n7805));
  orx   g06977(.a(n7805), .b(n7804), .O(n7806));
  andx  g06978(.a(n7806), .b(n7792), .O(n7807));
  andx  g06979(.a(n7807), .b(n7784), .O(n7808));
  orx   g06980(.a(n7618), .b(n7616), .O(n7809));
  orx   g06981(.a(n7619), .b(n7635), .O(n7810));
  andx  g06982(.a(n7810), .b(n7809), .O(n7811));
  orx   g06983(.a(n7811), .b(n7632), .O(n7812));
  andx  g06984(.a(n7619), .b(n7635), .O(n7813));
  andx  g06985(.a(n7618), .b(n7616), .O(n7814));
  orx   g06986(.a(n7814), .b(n7813), .O(n7815));
  orx   g06987(.a(n7815), .b(n7340), .O(n7816));
  andx  g06988(.a(n7816), .b(n7812), .O(n7817));
  andx  g06989(.a(n7817), .b(n7808), .O(n7818));
  orx   g06990(.a(n7624), .b(n7622), .O(n7819));
  andx  g06991(.a(n7625), .b(n7819), .O(n7821));
  orx   g06992(.a(n7821), .b(n7629), .O(n7822));
  andx  g06993(.a(n7625), .b(n7639), .O(n7823));
  orx   g06994(.a(n7624), .b(n7823), .O(n7825));
  orx   g06995(.a(n7825), .b(n7331), .O(n7826));
  andx  g06996(.a(n7826), .b(n7822), .O(n7827));
  andx  g06997(.a(n7827), .b(n7818), .O(n7828));
  orx   g06998(.a(n7641), .b(n7315), .O(n7829));
  andx  g06999(.a(n7308), .b(n7293), .O(n7831));
  orx   g07000(.a(n7831), .b(n7259), .O(n7832));
  orx   g07001(.a(n7640), .b(n7832), .O(n7833));
  andx  g07002(.a(n7833), .b(n7829), .O(n7834));
  andx  g07003(.a(n7834), .b(n7828), .O(n7835));
  andx  g07004(.a(n7259), .b(n7290), .O(n7836));
  invx  g07005(.a(n7836), .O(n7837));
  orx   g07006(.a(n7259), .b(n7290), .O(n7838));
  andx  g07007(.a(n7838), .b(n7740), .O(n7839));
  andx  g07008(.a(n7839), .b(n7837), .O(n7840));
  orx   g07009(.a(n7840), .b(n7646), .O(n7841));
  andx  g07010(.a(n7841), .b(n7835), .O(n7842));
  orx   g07011(.a(n7261), .b(n7768), .O(n7843));
  orx   g07012(.a(n7843), .b(n7646), .O(n7844));
  orx   g07013(.a(n7306), .b(n6933), .O(n7845));
  orx   g07014(.a(n7742), .b(n6933), .O(n7846));
  andx  g07015(.a(n7846), .b(n7845), .O(n7847));
  andx  g07016(.a(n7847), .b(n7844), .O(n7848));
  andx  g07017(.a(n7848), .b(n7842), .O(n7849));
  andx  g07018(.a(n7849), .b(n7775), .O(n7850));
  invx  g07019(.a(n6572), .O(n7851));
  orx   g07020(.a(n6591), .b(n6573), .O(n7852));
  orx   g07021(.a(n6587), .b(n6239), .O(n7853));
  andx  g07022(.a(n7853), .b(n7852), .O(n7854));
  orx   g07023(.a(n7854), .b(n7851), .O(n7855));
  andx  g07024(.a(n7855), .b(n6594), .O(n7856));
  andx  g07025(.a(n7773), .b(n7270), .O(n7857));
  orx   g07026(.a(n7857), .b(n7273), .O(n7858));
  invx  g07027(.a(n7858), .O(n7859));
  orx   g07028(.a(n7859), .b(n7856), .O(n7860));
  andx  g07029(.a(n7854), .b(n7851), .O(n7861));
  orx   g07030(.a(n7276), .b(n7861), .O(n7862));
  orx   g07031(.a(n7858), .b(n7862), .O(n7863));
  andx  g07032(.a(n7863), .b(n7860), .O(n7864));
  andx  g07033(.a(n7864), .b(n7850), .O(n7865));
  andx  g07034(.a(n7858), .b(n6594), .O(n7866));
  orx   g07035(.a(n7866), .b(n7278), .O(n7867));
  andx  g07036(.a(n7867), .b(n7286), .O(n7868));
  invx  g07037(.a(n7868), .O(n7869));
  orx   g07038(.a(n7867), .b(n7286), .O(n7870));
  andx  g07039(.a(n7870), .b(n7869), .O(n7871));
  invx  g07040(.a(n7871), .O(n7872));
  andx  g07041(.a(n7872), .b(n7865), .O(n7873));
  orx   g07042(.a(n5777), .b(n7737), .O(n7874));
  orx   g07043(.a(n7874), .b(n7868), .O(n7875));
  orx   g07044(.a(n7738), .b(n5397), .O(n7876));
  orx   g07045(.a(n7869), .b(n5397), .O(n7877));
  andx  g07046(.a(n7877), .b(n7876), .O(n7878));
  andx  g07047(.a(n7878), .b(n7875), .O(n7879));
  andx  g07048(.a(n7879), .b(n7873), .O(n7880));
  andx  g07049(.a(n7880), .b(n7763), .O(n7881));
  andx  g07050(.a(n7761), .b(n5390), .O(n7882));
  orx   g07051(.a(n7882), .b(n5389), .O(n7883));
  invx  g07052(.a(n5781), .O(n7884));
  orx   g07053(.a(n7884), .b(n5077), .O(n7885));
  andx  g07054(.a(n7885), .b(n7883), .O(n7886));
  invx  g07055(.a(n7886), .O(n7887));
  orx   g07056(.a(n7885), .b(n7883), .O(n7888));
  andx  g07057(.a(n7888), .b(n7887), .O(n7889));
  andx  g07058(.a(n7889), .b(n7881), .O(n7890));
  andx  g07059(.a(n7883), .b(n5781), .O(n7891));
  orx   g07060(.a(n7891), .b(n5079), .O(n7892));
  andx  g07061(.a(n7892), .b(n5866), .O(n7893));
  invx  g07062(.a(n7893), .O(n7894));
  orx   g07063(.a(n7892), .b(n5866), .O(n7895));
  andx  g07064(.a(n7895), .b(n7894), .O(n7896));
  invx  g07065(.a(n7896), .O(n7897));
  andx  g07066(.a(n7897), .b(n7890), .O(n7898));
  invx  g07067(.a(n7898), .O(n7899));
  andx  g07068(.a(n7899), .b(n7732), .O(n7900));
  andx  g07069(.a(n7898), .b(n7731), .O(n7901));
  orx   g07070(.a(n7901), .b(n7900), .O(n7902));
  andx  g07071(.a(n7902), .b(n1790), .O(n7903));
  orx   g07072(.a(n7871), .b(n7865), .O(n7904));
  invx  g07073(.a(n7904), .O(n7905));
  andx  g07074(.a(n7871), .b(n7865), .O(n7906));
  orx   g07075(.a(n7906), .b(n7905), .O(n7907));
  andx  g07076(.a(n7907), .b(n3210), .O(n7908));
  invx  g07077(.a(n7908), .O(n7909));
  invx  g07078(.a(n7818), .O(n7910));
  orx   g07079(.a(n7827), .b(n7910), .O(n7911));
  andx  g07080(.a(n7825), .b(n7331), .O(n7912));
  andx  g07081(.a(n7821), .b(n7629), .O(n7913));
  orx   g07082(.a(n7913), .b(n7912), .O(n7914));
  orx   g07083(.a(n7914), .b(n7818), .O(n7915));
  andx  g07084(.a(n7915), .b(n7911), .O(n7916));
  orx   g07085(.a(n7916), .b(n3418), .O(n7917));
  invx  g07086(.a(n7808), .O(n7918));
  andx  g07087(.a(n7817), .b(n7918), .O(n7919));
  andx  g07088(.a(n7815), .b(n7340), .O(n7920));
  andx  g07089(.a(n7811), .b(n7632), .O(n7921));
  orx   g07090(.a(n7921), .b(n7920), .O(n7922));
  andx  g07091(.a(n7922), .b(n7808), .O(n7923));
  orx   g07092(.a(n7923), .b(n7919), .O(n7924));
  andx  g07093(.a(n7782), .b(n7534), .O(n7925));
  andx  g07094(.a(n7778), .b(n7611), .O(n7926));
  orx   g07095(.a(n7926), .b(n7925), .O(n7927));
  andx  g07096(.a(n7807), .b(n7927), .O(n7928));
  invx  g07097(.a(n7807), .O(n7929));
  andx  g07098(.a(n7929), .b(n7784), .O(n7930));
  orx   g07099(.a(n7930), .b(n7928), .O(n7931));
  andx  g07100(.a(n7931), .b(n3171), .O(n7932));
  andx  g07101(.a(n7791), .b(n3645), .O(n7933));
  invx  g07102(.a(n7805), .O(n7934));
  andx  g07103(.a(n7934), .b(n7803), .O(n7935));
  andx  g07104(.a(n7935), .b(n7792), .O(n7936));
  andx  g07105(.a(n7806), .b(n7791), .O(n7937));
  orx   g07106(.a(n7937), .b(n7936), .O(n7938));
  andx  g07107(.a(n7938), .b(n3413), .O(n7939));
  orx   g07108(.a(n7939), .b(n7933), .O(n7940));
  andx  g07109(.a(n7939), .b(n7933), .O(n7941));
  invx  g07110(.a(n7941), .O(n7942));
  andx  g07111(.a(n7942), .b(n7940), .O(n7943));
  andx  g07112(.a(n7943), .b(n7932), .O(n7944));
  andx  g07113(.a(n7791), .b(n3413), .O(n7945));
  andx  g07114(.a(n7938), .b(n3171), .O(n7946));
  andx  g07115(.a(n7946), .b(n7945), .O(n7947));
  andx  g07116(.a(n7947), .b(n7932), .O(n7948));
  andx  g07117(.a(n7947), .b(n7943), .O(n7949));
  orx   g07118(.a(n7949), .b(n7948), .O(n7950));
  orx   g07119(.a(n7950), .b(n7944), .O(n7951));
  andx  g07120(.a(n7951), .b(n7924), .O(n7952));
  andx  g07121(.a(n7924), .b(n3171), .O(n7953));
  orx   g07122(.a(n7953), .b(n7951), .O(n7954));
  andx  g07123(.a(n7931), .b(n3413), .O(n7955));
  andx  g07124(.a(n7955), .b(n7942), .O(n7956));
  orx   g07125(.a(n7929), .b(n7784), .O(n7957));
  orx   g07126(.a(n7807), .b(n7927), .O(n7958));
  andx  g07127(.a(n7958), .b(n7957), .O(n7959));
  orx   g07128(.a(n7959), .b(n4989), .O(n7960));
  andx  g07129(.a(n7960), .b(n7941), .O(n7961));
  orx   g07130(.a(n7961), .b(n7956), .O(n7962));
  andx  g07131(.a(n7791), .b(n3721), .O(n7963));
  invx  g07132(.a(n7963), .O(n7964));
  andx  g07133(.a(n7938), .b(n3645), .O(n7965));
  orx   g07134(.a(n7965), .b(n7964), .O(n7966));
  orx   g07135(.a(n7806), .b(n7791), .O(n7967));
  orx   g07136(.a(n7935), .b(n7792), .O(n7968));
  andx  g07137(.a(n7968), .b(n7967), .O(n7969));
  orx   g07138(.a(n7969), .b(n4509), .O(n7970));
  orx   g07139(.a(n7970), .b(n7963), .O(n7971));
  andx  g07140(.a(n7971), .b(n7966), .O(n7972));
  orx   g07141(.a(n7972), .b(n7962), .O(n7973));
  invx  g07142(.a(n7973), .O(n7974));
  andx  g07143(.a(n7972), .b(n7962), .O(n7975));
  orx   g07144(.a(n7975), .b(n7974), .O(n7976));
  andx  g07145(.a(n7976), .b(n7954), .O(n7977));
  orx   g07146(.a(n7977), .b(n7952), .O(n7978));
  orx   g07147(.a(n7978), .b(n7917), .O(n7979));
  andx  g07148(.a(n7914), .b(n7818), .O(n7980));
  andx  g07149(.a(n7827), .b(n7910), .O(n7981));
  orx   g07150(.a(n7981), .b(n7980), .O(n7982));
  andx  g07151(.a(n7982), .b(n3171), .O(n7983));
  invx  g07152(.a(n7952), .O(n7984));
  invx  g07153(.a(n7944), .O(n7985));
  invx  g07154(.a(n7948), .O(n7986));
  invx  g07155(.a(n7940), .O(n7987));
  orx   g07156(.a(n7941), .b(n7987), .O(n7988));
  invx  g07157(.a(n7947), .O(n7989));
  orx   g07158(.a(n7989), .b(n7988), .O(n7990));
  andx  g07159(.a(n7990), .b(n7986), .O(n7991));
  andx  g07160(.a(n7991), .b(n7985), .O(n7992));
  invx  g07161(.a(n7953), .O(n7993));
  andx  g07162(.a(n7993), .b(n7992), .O(n7994));
  invx  g07163(.a(n7975), .O(n7995));
  andx  g07164(.a(n7995), .b(n7973), .O(n7996));
  orx   g07165(.a(n7996), .b(n7994), .O(n7997));
  andx  g07166(.a(n7997), .b(n7984), .O(n7998));
  orx   g07167(.a(n7998), .b(n7983), .O(n7999));
  andx  g07168(.a(n7999), .b(n7979), .O(n8000));
  andx  g07169(.a(n7955), .b(n7941), .O(n8001));
  invx  g07170(.a(n8001), .O(n8002));
  orx   g07171(.a(n7972), .b(n7960), .O(n8003));
  orx   g07172(.a(n7972), .b(n7942), .O(n8004));
  andx  g07173(.a(n8004), .b(n8003), .O(n8005));
  andx  g07174(.a(n8005), .b(n8002), .O(n8006));
  orx   g07175(.a(n7922), .b(n7808), .O(n8007));
  orx   g07176(.a(n7817), .b(n7918), .O(n8008));
  andx  g07177(.a(n8008), .b(n8007), .O(n8009));
  orx   g07178(.a(n8009), .b(n4989), .O(n8010));
  andx  g07179(.a(n8010), .b(n8006), .O(n8011));
  andx  g07180(.a(n7970), .b(n7963), .O(n8012));
  andx  g07181(.a(n7965), .b(n7964), .O(n8013));
  orx   g07182(.a(n8013), .b(n8012), .O(n8014));
  andx  g07183(.a(n8014), .b(n7955), .O(n8015));
  andx  g07184(.a(n8014), .b(n7941), .O(n8016));
  orx   g07185(.a(n8016), .b(n8015), .O(n8017));
  orx   g07186(.a(n8017), .b(n8001), .O(n8018));
  andx  g07187(.a(n8018), .b(n7924), .O(n8019));
  orx   g07188(.a(n8019), .b(n8011), .O(n8020));
  andx  g07189(.a(n7965), .b(n7963), .O(n8021));
  orx   g07190(.a(n7959), .b(n4509), .O(n8022));
  orx   g07191(.a(n8022), .b(n8021), .O(n8023));
  invx  g07192(.a(n8021), .O(n8024));
  andx  g07193(.a(n7931), .b(n3645), .O(n8025));
  orx   g07194(.a(n8025), .b(n8024), .O(n8026));
  andx  g07195(.a(n8026), .b(n8023), .O(n8027));
  andx  g07196(.a(n7791), .b(n4063), .O(n8028));
  orx   g07197(.a(n7969), .b(n6829), .O(n8029));
  andx  g07198(.a(n8029), .b(n8028), .O(n8030));
  invx  g07199(.a(n8028), .O(n8031));
  andx  g07200(.a(n7938), .b(n3721), .O(n8032));
  andx  g07201(.a(n8032), .b(n8031), .O(n8033));
  orx   g07202(.a(n8033), .b(n8030), .O(n8034));
  andx  g07203(.a(n8034), .b(n8027), .O(n8035));
  andx  g07204(.a(n8025), .b(n8024), .O(n8036));
  andx  g07205(.a(n8022), .b(n8021), .O(n8037));
  orx   g07206(.a(n8037), .b(n8036), .O(n8038));
  orx   g07207(.a(n8032), .b(n8031), .O(n8039));
  orx   g07208(.a(n8029), .b(n8028), .O(n8040));
  andx  g07209(.a(n8040), .b(n8039), .O(n8041));
  andx  g07210(.a(n8041), .b(n8038), .O(n8042));
  orx   g07211(.a(n8042), .b(n8035), .O(n8043));
  andx  g07212(.a(n8043), .b(n8020), .O(n8044));
  invx  g07213(.a(n8044), .O(n8045));
  orx   g07214(.a(n8043), .b(n8020), .O(n8046));
  andx  g07215(.a(n8046), .b(n8045), .O(n8047));
  orx   g07216(.a(n8047), .b(n8000), .O(n8048));
  andx  g07217(.a(n7998), .b(n7983), .O(n8049));
  andx  g07218(.a(n7978), .b(n7917), .O(n8050));
  orx   g07219(.a(n8050), .b(n8049), .O(n8051));
  invx  g07220(.a(n8046), .O(n8052));
  orx   g07221(.a(n8052), .b(n8044), .O(n8053));
  orx   g07222(.a(n8053), .b(n8051), .O(n8054));
  andx  g07223(.a(n8054), .b(n8048), .O(n8055));
  invx  g07224(.a(n7828), .O(n8056));
  andx  g07225(.a(n7834), .b(n8056), .O(n8057));
  andx  g07226(.a(n7640), .b(n7832), .O(n8058));
  andx  g07227(.a(n7641), .b(n7315), .O(n8059));
  orx   g07228(.a(n8059), .b(n8058), .O(n8060));
  andx  g07229(.a(n8060), .b(n7828), .O(n8061));
  orx   g07230(.a(n8061), .b(n8057), .O(n8062));
  andx  g07231(.a(n8062), .b(n3429), .O(n8063));
  andx  g07232(.a(n7982), .b(n3429), .O(n8064));
  andx  g07233(.a(n7931), .b(n3429), .O(n8065));
  orx   g07234(.a(n7946), .b(n7945), .O(n8066));
  andx  g07235(.a(n8066), .b(n7989), .O(n8067));
  andx  g07236(.a(n8067), .b(n8065), .O(n8068));
  andx  g07237(.a(n7791), .b(n3171), .O(n8069));
  andx  g07238(.a(n7938), .b(n3429), .O(n8070));
  andx  g07239(.a(n8070), .b(n8069), .O(n8071));
  andx  g07240(.a(n8071), .b(n8065), .O(n8072));
  andx  g07241(.a(n8071), .b(n8067), .O(n8073));
  orx   g07242(.a(n8073), .b(n8072), .O(n8074));
  orx   g07243(.a(n8074), .b(n8068), .O(n8075));
  andx  g07244(.a(n8075), .b(n7924), .O(n8076));
  andx  g07245(.a(n7989), .b(n7932), .O(n8077));
  invx  g07246(.a(n8077), .O(n8078));
  orx   g07247(.a(n7989), .b(n7932), .O(n8079));
  andx  g07248(.a(n8079), .b(n8078), .O(n8080));
  andx  g07249(.a(n8080), .b(n7943), .O(n8081));
  orx   g07250(.a(n8080), .b(n7943), .O(n8082));
  invx  g07251(.a(n8082), .O(n8083));
  orx   g07252(.a(n8083), .b(n8081), .O(n8084));
  andx  g07253(.a(n7924), .b(n3429), .O(n8085));
  orx   g07254(.a(n8085), .b(n8075), .O(n8086));
  andx  g07255(.a(n8086), .b(n8084), .O(n8087));
  orx   g07256(.a(n8087), .b(n8076), .O(n8088));
  andx  g07257(.a(n8088), .b(n8064), .O(n8089));
  orx   g07258(.a(n7994), .b(n7952), .O(n8090));
  andx  g07259(.a(n8090), .b(n7976), .O(n8091));
  orx   g07260(.a(n8090), .b(n7976), .O(n8092));
  invx  g07261(.a(n8092), .O(n8093));
  orx   g07262(.a(n8093), .b(n8091), .O(n8094));
  orx   g07263(.a(n8088), .b(n8064), .O(n8095));
  andx  g07264(.a(n8095), .b(n8094), .O(n8096));
  orx   g07265(.a(n8096), .b(n8089), .O(n8097));
  andx  g07266(.a(n8097), .b(n8063), .O(n8098));
  invx  g07267(.a(n8063), .O(n8099));
  invx  g07268(.a(n8089), .O(n8100));
  invx  g07269(.a(n8091), .O(n8101));
  andx  g07270(.a(n8092), .b(n8101), .O(n8102));
  invx  g07271(.a(n8064), .O(n8103));
  invx  g07272(.a(n8076), .O(n8104));
  invx  g07273(.a(n8081), .O(n8105));
  andx  g07274(.a(n8082), .b(n8105), .O(n8106));
  invx  g07275(.a(n8086), .O(n8107));
  orx   g07276(.a(n8107), .b(n8106), .O(n8108));
  andx  g07277(.a(n8108), .b(n8104), .O(n8109));
  andx  g07278(.a(n8109), .b(n8103), .O(n8110));
  orx   g07279(.a(n8110), .b(n8102), .O(n8111));
  andx  g07280(.a(n8111), .b(n8100), .O(n8112));
  andx  g07281(.a(n8112), .b(n8099), .O(n8113));
  orx   g07282(.a(n8113), .b(n8098), .O(n8114));
  andx  g07283(.a(n8114), .b(n8055), .O(n8115));
  andx  g07284(.a(n8053), .b(n8051), .O(n8116));
  andx  g07285(.a(n8047), .b(n8000), .O(n8117));
  orx   g07286(.a(n8117), .b(n8116), .O(n8118));
  orx   g07287(.a(n8112), .b(n8099), .O(n8119));
  orx   g07288(.a(n8097), .b(n8063), .O(n8120));
  andx  g07289(.a(n8120), .b(n8119), .O(n8121));
  andx  g07290(.a(n8121), .b(n8118), .O(n8122));
  orx   g07291(.a(n8122), .b(n8115), .O(n8123));
  invx  g07292(.a(n7835), .O(n8124));
  andx  g07293(.a(n7841), .b(n8124), .O(n8125));
  andx  g07294(.a(n7310), .b(n6942), .O(n8126));
  orx   g07295(.a(n8126), .b(n7644), .O(n8127));
  orx   g07296(.a(n8127), .b(n7836), .O(n8128));
  andx  g07297(.a(n8128), .b(n7742), .O(n8129));
  andx  g07298(.a(n8129), .b(n7835), .O(n8130));
  orx   g07299(.a(n8130), .b(n8125), .O(n8131));
  andx  g07300(.a(n8131), .b(n3180), .O(n8132));
  andx  g07301(.a(n8132), .b(n8123), .O(n8133));
  invx  g07302(.a(n8133), .O(n8134));
  orx   g07303(.a(n8121), .b(n8118), .O(n8135));
  orx   g07304(.a(n8114), .b(n8055), .O(n8136));
  andx  g07305(.a(n8136), .b(n8135), .O(n8137));
  orx   g07306(.a(n8088), .b(n8103), .O(n8138));
  orx   g07307(.a(n8109), .b(n8064), .O(n8139));
  andx  g07308(.a(n8139), .b(n8138), .O(n8140));
  orx   g07309(.a(n8140), .b(n8102), .O(n8141));
  andx  g07310(.a(n8109), .b(n8064), .O(n8142));
  andx  g07311(.a(n8088), .b(n8103), .O(n8143));
  orx   g07312(.a(n8143), .b(n8142), .O(n8144));
  orx   g07313(.a(n8144), .b(n8094), .O(n8145));
  andx  g07314(.a(n8145), .b(n8141), .O(n8146));
  andx  g07315(.a(n7982), .b(n3180), .O(n8147));
  andx  g07316(.a(n7931), .b(n3180), .O(n8148));
  invx  g07317(.a(n8070), .O(n8149));
  andx  g07318(.a(n8149), .b(n8069), .O(n8150));
  invx  g07319(.a(n8069), .O(n8151));
  andx  g07320(.a(n8070), .b(n8151), .O(n8152));
  orx   g07321(.a(n8152), .b(n8150), .O(n8153));
  andx  g07322(.a(n8153), .b(n8148), .O(n8154));
  andx  g07323(.a(n7791), .b(n3429), .O(n8155));
  andx  g07324(.a(n7938), .b(n3180), .O(n8156));
  andx  g07325(.a(n8156), .b(n8155), .O(n8157));
  andx  g07326(.a(n8157), .b(n8148), .O(n8158));
  andx  g07327(.a(n8157), .b(n8153), .O(n8159));
  orx   g07328(.a(n8159), .b(n8158), .O(n8160));
  orx   g07329(.a(n8160), .b(n8154), .O(n8161));
  andx  g07330(.a(n8161), .b(n7924), .O(n8162));
  invx  g07331(.a(n8162), .O(n8163));
  invx  g07332(.a(n8067), .O(n8164));
  invx  g07333(.a(n8071), .O(n8165));
  andx  g07334(.a(n8165), .b(n8065), .O(n8166));
  invx  g07335(.a(n8065), .O(n8167));
  andx  g07336(.a(n8071), .b(n8167), .O(n8168));
  orx   g07337(.a(n8168), .b(n8166), .O(n8169));
  orx   g07338(.a(n8169), .b(n8164), .O(n8170));
  andx  g07339(.a(n8169), .b(n8164), .O(n8171));
  invx  g07340(.a(n8171), .O(n8172));
  andx  g07341(.a(n8172), .b(n8170), .O(n8173));
  andx  g07342(.a(n7924), .b(n3180), .O(n8174));
  orx   g07343(.a(n8174), .b(n8161), .O(n8175));
  invx  g07344(.a(n8175), .O(n8176));
  orx   g07345(.a(n8176), .b(n8173), .O(n8177));
  andx  g07346(.a(n8177), .b(n8163), .O(n8178));
  invx  g07347(.a(n8178), .O(n8179));
  andx  g07348(.a(n8179), .b(n8147), .O(n8180));
  andx  g07349(.a(n8086), .b(n8104), .O(n8181));
  orx   g07350(.a(n8181), .b(n8106), .O(n8182));
  invx  g07351(.a(n8182), .O(n8183));
  andx  g07352(.a(n8181), .b(n8106), .O(n8184));
  orx   g07353(.a(n8184), .b(n8183), .O(n8185));
  invx  g07354(.a(n8147), .O(n8186));
  andx  g07355(.a(n8178), .b(n8186), .O(n8187));
  invx  g07356(.a(n8187), .O(n8188));
  andx  g07357(.a(n8188), .b(n8185), .O(n8189));
  orx   g07358(.a(n8189), .b(n8180), .O(n8190));
  andx  g07359(.a(n8190), .b(n8146), .O(n8191));
  invx  g07360(.a(n8191), .O(n8192));
  andx  g07361(.a(n8144), .b(n8094), .O(n8193));
  andx  g07362(.a(n8140), .b(n8102), .O(n8194));
  orx   g07363(.a(n8194), .b(n8193), .O(n8195));
  invx  g07364(.a(n8180), .O(n8196));
  invx  g07365(.a(n8184), .O(n8197));
  andx  g07366(.a(n8197), .b(n8182), .O(n8198));
  orx   g07367(.a(n8187), .b(n8198), .O(n8199));
  andx  g07368(.a(n8199), .b(n8196), .O(n8200));
  andx  g07369(.a(n8200), .b(n8195), .O(n8201));
  andx  g07370(.a(n8062), .b(n3180), .O(n8202));
  invx  g07371(.a(n8202), .O(n8203));
  orx   g07372(.a(n8203), .b(n8201), .O(n8204));
  andx  g07373(.a(n8204), .b(n8192), .O(n8205));
  orx   g07374(.a(n8205), .b(n8137), .O(n8206));
  invx  g07375(.a(n8132), .O(n8207));
  orx   g07376(.a(n8205), .b(n8207), .O(n8208));
  andx  g07377(.a(n8208), .b(n8206), .O(n8209));
  andx  g07378(.a(n8209), .b(n8134), .O(n8210));
  invx  g07379(.a(n7842), .O(n8211));
  andx  g07380(.a(n7306), .b(n6933), .O(n8212));
  andx  g07381(.a(n8212), .b(n7742), .O(n8213));
  andx  g07382(.a(n7261), .b(n7768), .O(n8214));
  andx  g07383(.a(n7646), .b(n7768), .O(n8215));
  orx   g07384(.a(n8215), .b(n8214), .O(n8216));
  orx   g07385(.a(n8216), .b(n8213), .O(n8217));
  orx   g07386(.a(n8217), .b(n8211), .O(n8218));
  orx   g07387(.a(n7848), .b(n7842), .O(n8219));
  andx  g07388(.a(n8219), .b(n8218), .O(n8220));
  andx  g07389(.a(n8220), .b(n3180), .O(n8221));
  andx  g07390(.a(n8221), .b(n8210), .O(n8222));
  orx   g07391(.a(n8190), .b(n8146), .O(n8223));
  andx  g07392(.a(n8202), .b(n8223), .O(n8224));
  orx   g07393(.a(n8224), .b(n8191), .O(n8225));
  andx  g07394(.a(n8225), .b(n8123), .O(n8226));
  andx  g07395(.a(n8225), .b(n8132), .O(n8227));
  orx   g07396(.a(n8227), .b(n8226), .O(n8228));
  orx   g07397(.a(n8228), .b(n8133), .O(n8229));
  invx  g07398(.a(n8221), .O(n8230));
  andx  g07399(.a(n8230), .b(n8229), .O(n8231));
  orx   g07400(.a(n8231), .b(n8222), .O(n8232));
  andx  g07401(.a(n7982), .b(n3413), .O(n8233));
  invx  g07402(.a(n8019), .O(n8234));
  orx   g07403(.a(n8041), .b(n8038), .O(n8235));
  orx   g07404(.a(n8034), .b(n8027), .O(n8236));
  andx  g07405(.a(n8236), .b(n8235), .O(n8237));
  orx   g07406(.a(n8237), .b(n8011), .O(n8238));
  andx  g07407(.a(n8238), .b(n8234), .O(n8239));
  andx  g07408(.a(n8239), .b(n8233), .O(n8240));
  orx   g07409(.a(n7916), .b(n4989), .O(n8241));
  andx  g07410(.a(n7924), .b(n3413), .O(n8242));
  orx   g07411(.a(n8242), .b(n8018), .O(n8243));
  andx  g07412(.a(n8043), .b(n8243), .O(n8244));
  orx   g07413(.a(n8244), .b(n8019), .O(n8245));
  andx  g07414(.a(n8245), .b(n8241), .O(n8246));
  orx   g07415(.a(n8246), .b(n8240), .O(n8247));
  andx  g07416(.a(n8025), .b(n8021), .O(n8248));
  invx  g07417(.a(n8248), .O(n8249));
  orx   g07418(.a(n8041), .b(n8022), .O(n8250));
  orx   g07419(.a(n8041), .b(n8024), .O(n8251));
  andx  g07420(.a(n8251), .b(n8250), .O(n8252));
  andx  g07421(.a(n8252), .b(n8249), .O(n8253));
  orx   g07422(.a(n8009), .b(n4509), .O(n8254));
  andx  g07423(.a(n8254), .b(n8253), .O(n8255));
  andx  g07424(.a(n8034), .b(n8025), .O(n8256));
  andx  g07425(.a(n8034), .b(n8021), .O(n8257));
  orx   g07426(.a(n8257), .b(n8256), .O(n8258));
  orx   g07427(.a(n8258), .b(n8248), .O(n8259));
  andx  g07428(.a(n8259), .b(n7924), .O(n8260));
  orx   g07429(.a(n8260), .b(n8255), .O(n8261));
  andx  g07430(.a(n8032), .b(n8028), .O(n8262));
  orx   g07431(.a(n7959), .b(n6829), .O(n8263));
  orx   g07432(.a(n8263), .b(n8262), .O(n8264));
  invx  g07433(.a(n8262), .O(n8265));
  andx  g07434(.a(n7931), .b(n3721), .O(n8266));
  orx   g07435(.a(n8266), .b(n8265), .O(n8267));
  andx  g07436(.a(n8267), .b(n8264), .O(n8268));
  andx  g07437(.a(n7791), .b(n4114), .O(n8269));
  orx   g07438(.a(n7969), .b(n4062), .O(n8270));
  andx  g07439(.a(n8270), .b(n8269), .O(n8271));
  invx  g07440(.a(n8269), .O(n8272));
  andx  g07441(.a(n7938), .b(n4063), .O(n8273));
  andx  g07442(.a(n8273), .b(n8272), .O(n8274));
  orx   g07443(.a(n8274), .b(n8271), .O(n8275));
  andx  g07444(.a(n8275), .b(n8268), .O(n8276));
  andx  g07445(.a(n8266), .b(n8265), .O(n8277));
  andx  g07446(.a(n8263), .b(n8262), .O(n8278));
  orx   g07447(.a(n8278), .b(n8277), .O(n8279));
  orx   g07448(.a(n8273), .b(n8272), .O(n8280));
  orx   g07449(.a(n8270), .b(n8269), .O(n8281));
  andx  g07450(.a(n8281), .b(n8280), .O(n8282));
  andx  g07451(.a(n8282), .b(n8279), .O(n8283));
  orx   g07452(.a(n8283), .b(n8276), .O(n8284));
  andx  g07453(.a(n8284), .b(n8261), .O(n8285));
  orx   g07454(.a(n8284), .b(n8261), .O(n8286));
  invx  g07455(.a(n8286), .O(n8287));
  orx   g07456(.a(n8287), .b(n8285), .O(n8288));
  andx  g07457(.a(n8288), .b(n8247), .O(n8289));
  orx   g07458(.a(n8245), .b(n8241), .O(n8290));
  orx   g07459(.a(n8239), .b(n8233), .O(n8291));
  andx  g07460(.a(n8291), .b(n8290), .O(n8292));
  invx  g07461(.a(n8285), .O(n8293));
  andx  g07462(.a(n8286), .b(n8293), .O(n8294));
  andx  g07463(.a(n8294), .b(n8292), .O(n8295));
  orx   g07464(.a(n8295), .b(n8289), .O(n8296));
  orx   g07465(.a(n8060), .b(n7828), .O(n8297));
  orx   g07466(.a(n7834), .b(n8056), .O(n8298));
  andx  g07467(.a(n8298), .b(n8297), .O(n8299));
  orx   g07468(.a(n8299), .b(n3418), .O(n8300));
  andx  g07469(.a(n7978), .b(n7983), .O(n8301));
  orx   g07470(.a(n7978), .b(n7983), .O(n8302));
  andx  g07471(.a(n8302), .b(n8053), .O(n8303));
  orx   g07472(.a(n8303), .b(n8301), .O(n8304));
  andx  g07473(.a(n8304), .b(n8300), .O(n8305));
  andx  g07474(.a(n8062), .b(n3171), .O(n8306));
  invx  g07475(.a(n8301), .O(n8307));
  andx  g07476(.a(n7998), .b(n7917), .O(n8308));
  orx   g07477(.a(n8308), .b(n8047), .O(n8309));
  andx  g07478(.a(n8309), .b(n8307), .O(n8310));
  andx  g07479(.a(n8310), .b(n8306), .O(n8311));
  orx   g07480(.a(n8311), .b(n8305), .O(n8312));
  andx  g07481(.a(n8312), .b(n8296), .O(n8313));
  orx   g07482(.a(n8312), .b(n8296), .O(n8315));
  andx  g07483(.a(n8131), .b(n3429), .O(n8317));
  invx  g07484(.a(n8317), .O(n8318));
  andx  g07485(.a(n8097), .b(n8055), .O(n8319));
  orx   g07486(.a(n8097), .b(n8055), .O(n8320));
  andx  g07487(.a(n8320), .b(n8063), .O(n8321));
  orx   g07488(.a(n8321), .b(n8319), .O(n8322));
  andx  g07489(.a(n8322), .b(n8318), .O(n8323));
  invx  g07490(.a(n8319), .O(n8324));
  andx  g07491(.a(n8112), .b(n8118), .O(n8325));
  orx   g07492(.a(n8325), .b(n8099), .O(n8326));
  andx  g07493(.a(n8326), .b(n8324), .O(n8327));
  andx  g07494(.a(n8327), .b(n8317), .O(n8328));
  orx   g07495(.a(n8328), .b(n8323), .O(n8329));
  andx  g07496(.a(n8329), .b(n8668), .O(n8330));
  orx   g07497(.a(n8327), .b(n8317), .O(n8332));
  orx   g07498(.a(n8322), .b(n8318), .O(n8333));
  andx  g07499(.a(n8333), .b(n8332), .O(n8334));
  andx  g07500(.a(n8334), .b(n8663), .O(n8335));
  orx   g07501(.a(n8335), .b(n8330), .O(n8336));
  andx  g07502(.a(n8336), .b(n8232), .O(n8337));
  orx   g07503(.a(n8230), .b(n8229), .O(n8338));
  orx   g07504(.a(n8221), .b(n8210), .O(n8339));
  andx  g07505(.a(n8339), .b(n8338), .O(n8340));
  orx   g07506(.a(n8334), .b(n8663), .O(n8341));
  orx   g07507(.a(n8329), .b(n8668), .O(n8342));
  andx  g07508(.a(n8342), .b(n8341), .O(n8343));
  andx  g07509(.a(n8343), .b(n8340), .O(n8344));
  orx   g07510(.a(n8344), .b(n8337), .O(n8345));
  andx  g07511(.a(n7773), .b(n7772), .O(n8346));
  andx  g07512(.a(n7770), .b(n7765), .O(n8347));
  orx   g07513(.a(n8347), .b(n8346), .O(n8348));
  orx   g07514(.a(n8218), .b(n8348), .O(n8349));
  orx   g07515(.a(n7849), .b(n7775), .O(n8350));
  andx  g07516(.a(n8350), .b(n8349), .O(n8351));
  andx  g07517(.a(n8351), .b(n3284), .O(n8352));
  invx  g07518(.a(n8352), .O(n8353));
  andx  g07519(.a(n8225), .b(n8207), .O(n8361));
  andx  g07520(.a(n8205), .b(n8132), .O(n8362));
  orx   g07521(.a(n8362), .b(n8361), .O(n8363));
  andx  g07522(.a(n8363), .b(n8137), .O(n8364));
  orx   g07523(.a(n8205), .b(n8132), .O(n8366));
  orx   g07524(.a(n8225), .b(n8207), .O(n8367));
  andx  g07525(.a(n8367), .b(n8366), .O(n8368));
  andx  g07526(.a(n8368), .b(n8123), .O(n8369));
  orx   g07527(.a(n8369), .b(n8364), .O(n8370));
  andx  g07528(.a(n8202), .b(n8190), .O(n8371));
  andx  g07529(.a(n8203), .b(n8200), .O(n8372));
  orx   g07530(.a(n8372), .b(n8371), .O(n8373));
  andx  g07531(.a(n8373), .b(n8146), .O(n8374));
  orx   g07532(.a(n8203), .b(n8200), .O(n8375));
  orx   g07533(.a(n8202), .b(n8190), .O(n8376));
  andx  g07534(.a(n8376), .b(n8375), .O(n8377));
  andx  g07535(.a(n8377), .b(n8195), .O(n8378));
  orx   g07536(.a(n8378), .b(n8374), .O(n8379));
  andx  g07537(.a(n8131), .b(n3284), .O(n8380));
  andx  g07538(.a(n8380), .b(n8379), .O(n8381));
  andx  g07539(.a(n8178), .b(n8147), .O(n8382));
  invx  g07540(.a(n8382), .O(n8383));
  orx   g07541(.a(n8178), .b(n8147), .O(n8384));
  andx  g07542(.a(n8384), .b(n8383), .O(n8385));
  orx   g07543(.a(n8385), .b(n8198), .O(n8386));
  invx  g07544(.a(n8384), .O(n8387));
  orx   g07545(.a(n8387), .b(n8382), .O(n8388));
  orx   g07546(.a(n8388), .b(n8185), .O(n8389));
  andx  g07547(.a(n8389), .b(n8386), .O(n8390));
  andx  g07548(.a(n8175), .b(n8163), .O(n8391));
  orx   g07549(.a(n8391), .b(n8173), .O(n8392));
  invx  g07550(.a(n8392), .O(n8393));
  andx  g07551(.a(n8391), .b(n8173), .O(n8394));
  orx   g07552(.a(n8394), .b(n8393), .O(n8395));
  andx  g07553(.a(n7931), .b(n3284), .O(n8396));
  invx  g07554(.a(n8156), .O(n8397));
  andx  g07555(.a(n8397), .b(n8155), .O(n8398));
  invx  g07556(.a(n8155), .O(n8399));
  andx  g07557(.a(n8156), .b(n8399), .O(n8400));
  orx   g07558(.a(n8400), .b(n8398), .O(n8401));
  andx  g07559(.a(n8401), .b(n8396), .O(n8402));
  andx  g07560(.a(n7791), .b(n3180), .O(n8403));
  andx  g07561(.a(n7938), .b(n3284), .O(n8404));
  andx  g07562(.a(n8404), .b(n8403), .O(n8405));
  andx  g07563(.a(n8405), .b(n8396), .O(n8406));
  andx  g07564(.a(n8405), .b(n8401), .O(n8407));
  orx   g07565(.a(n8407), .b(n8406), .O(n8408));
  orx   g07566(.a(n8408), .b(n8402), .O(n8409));
  andx  g07567(.a(n8409), .b(n7924), .O(n8410));
  invx  g07568(.a(n8157), .O(n8411));
  andx  g07569(.a(n8411), .b(n8148), .O(n8412));
  invx  g07570(.a(n8412), .O(n8413));
  orx   g07571(.a(n8411), .b(n8148), .O(n8414));
  andx  g07572(.a(n8414), .b(n8413), .O(n8415));
  andx  g07573(.a(n8149), .b(n8151), .O(n8416));
  orx   g07574(.a(n8416), .b(n8071), .O(n8417));
  andx  g07575(.a(n8417), .b(n8415), .O(n8418));
  invx  g07576(.a(n8418), .O(n8419));
  orx   g07577(.a(n8417), .b(n8415), .O(n8420));
  andx  g07578(.a(n8420), .b(n8419), .O(n8421));
  andx  g07579(.a(n7924), .b(n3284), .O(n8422));
  orx   g07580(.a(n8422), .b(n8409), .O(n8423));
  andx  g07581(.a(n8423), .b(n8421), .O(n8424));
  orx   g07582(.a(n8424), .b(n8410), .O(n8425));
  andx  g07583(.a(n8425), .b(n8395), .O(n8426));
  andx  g07584(.a(n7982), .b(n3284), .O(n8427));
  orx   g07585(.a(n8425), .b(n8395), .O(n8428));
  andx  g07586(.a(n8428), .b(n8427), .O(n8429));
  orx   g07587(.a(n8429), .b(n8426), .O(n8430));
  andx  g07588(.a(n8430), .b(n8390), .O(n8431));
  orx   g07589(.a(n8430), .b(n8390), .O(n8432));
  andx  g07590(.a(n8062), .b(n3284), .O(n8433));
  andx  g07591(.a(n8433), .b(n8432), .O(n8434));
  orx   g07592(.a(n8434), .b(n8431), .O(n8435));
  andx  g07593(.a(n8435), .b(n8379), .O(n8436));
  andx  g07594(.a(n8435), .b(n8380), .O(n8437));
  orx   g07595(.a(n8437), .b(n8436), .O(n8438));
  orx   g07596(.a(n8438), .b(n8381), .O(n8439));
  andx  g07597(.a(n8439), .b(n8370), .O(n8440));
  orx   g07598(.a(n8439), .b(n8370), .O(n8441));
  andx  g07599(.a(n8220), .b(n3284), .O(n8442));
  andx  g07600(.a(n8442), .b(n8441), .O(n8443));
  orx   g07601(.a(n8443), .b(n8440), .O(n8444));
  andx  g07602(.a(n8444), .b(n8353), .O(n8445));
  invx  g07603(.a(n8440), .O(n8446));
  orx   g07604(.a(n8368), .b(n8123), .O(n8447));
  orx   g07605(.a(n8363), .b(n8137), .O(n8448));
  andx  g07606(.a(n8448), .b(n8447), .O(n8449));
  invx  g07607(.a(n8381), .O(n8450));
  orx   g07608(.a(n8377), .b(n8195), .O(n8451));
  orx   g07609(.a(n8373), .b(n8146), .O(n8452));
  andx  g07610(.a(n8452), .b(n8451), .O(n8453));
  invx  g07611(.a(n8431), .O(n8454));
  andx  g07612(.a(n8388), .b(n8185), .O(n8455));
  andx  g07613(.a(n8385), .b(n8198), .O(n8456));
  orx   g07614(.a(n8456), .b(n8455), .O(n8457));
  invx  g07615(.a(n8426), .O(n8458));
  invx  g07616(.a(n8427), .O(n8459));
  invx  g07617(.a(n8394), .O(n8460));
  andx  g07618(.a(n8460), .b(n8392), .O(n8461));
  invx  g07619(.a(n8425), .O(n8462));
  andx  g07620(.a(n8462), .b(n8461), .O(n8463));
  orx   g07621(.a(n8463), .b(n8459), .O(n8464));
  andx  g07622(.a(n8464), .b(n8458), .O(n8465));
  andx  g07623(.a(n8465), .b(n8457), .O(n8466));
  invx  g07624(.a(n8433), .O(n8467));
  orx   g07625(.a(n8467), .b(n8466), .O(n8468));
  andx  g07626(.a(n8468), .b(n8454), .O(n8469));
  orx   g07627(.a(n8469), .b(n8453), .O(n8470));
  invx  g07628(.a(n8380), .O(n8471));
  orx   g07629(.a(n8469), .b(n8471), .O(n8472));
  andx  g07630(.a(n8472), .b(n8470), .O(n8473));
  andx  g07631(.a(n8473), .b(n8450), .O(n8474));
  andx  g07632(.a(n8474), .b(n8449), .O(n8475));
  invx  g07633(.a(n8442), .O(n8476));
  orx   g07634(.a(n8476), .b(n8475), .O(n8477));
  andx  g07635(.a(n8477), .b(n8446), .O(n8478));
  andx  g07636(.a(n8478), .b(n8352), .O(n8479));
  orx   g07637(.a(n8479), .b(n8445), .O(n8480));
  andx  g07638(.a(n8480), .b(n8345), .O(n8481));
  orx   g07639(.a(n8343), .b(n8340), .O(n8482));
  orx   g07640(.a(n8336), .b(n8232), .O(n8483));
  andx  g07641(.a(n8483), .b(n8482), .O(n8484));
  orx   g07642(.a(n8478), .b(n8352), .O(n8485));
  orx   g07643(.a(n8444), .b(n8353), .O(n8486));
  andx  g07644(.a(n8486), .b(n8485), .O(n8487));
  andx  g07645(.a(n8487), .b(n8484), .O(n8488));
  orx   g07646(.a(n8488), .b(n8481), .O(n8489));
  orx   g07647(.a(n8476), .b(n8439), .O(n8490));
  orx   g07648(.a(n8442), .b(n8474), .O(n8491));
  andx  g07649(.a(n8491), .b(n8490), .O(n8492));
  orx   g07650(.a(n8492), .b(n8449), .O(n8493));
  andx  g07651(.a(n8442), .b(n8474), .O(n8494));
  andx  g07652(.a(n8476), .b(n8439), .O(n8495));
  orx   g07653(.a(n8495), .b(n8494), .O(n8496));
  orx   g07654(.a(n8496), .b(n8370), .O(n8497));
  andx  g07655(.a(n8497), .b(n8493), .O(n8498));
  orx   g07656(.a(n8435), .b(n8380), .O(n8506));
  andx  g07657(.a(n8506), .b(n8472), .O(n8507));
  andx  g07658(.a(n8507), .b(n8453), .O(n8508));
  andx  g07659(.a(n8469), .b(n8471), .O(n8510));
  orx   g07660(.a(n8510), .b(n8437), .O(n8511));
  andx  g07661(.a(n8511), .b(n8379), .O(n8512));
  orx   g07662(.a(n8512), .b(n8508), .O(n8513));
  andx  g07663(.a(n8467), .b(n8430), .O(n8514));
  andx  g07664(.a(n8433), .b(n8465), .O(n8515));
  orx   g07665(.a(n8515), .b(n8514), .O(n8516));
  andx  g07666(.a(n8516), .b(n8457), .O(n8517));
  orx   g07667(.a(n8433), .b(n8465), .O(n8518));
  orx   g07668(.a(n8467), .b(n8430), .O(n8519));
  andx  g07669(.a(n8519), .b(n8518), .O(n8520));
  andx  g07670(.a(n8520), .b(n8390), .O(n8521));
  orx   g07671(.a(n8521), .b(n8517), .O(n8522));
  andx  g07672(.a(n8459), .b(n8425), .O(n8523));
  andx  g07673(.a(n8427), .b(n8462), .O(n8524));
  orx   g07674(.a(n8524), .b(n8523), .O(n8525));
  andx  g07675(.a(n8525), .b(n8395), .O(n8526));
  invx  g07676(.a(n8526), .O(n8527));
  orx   g07677(.a(n8525), .b(n8395), .O(n8528));
  andx  g07678(.a(n8528), .b(n8527), .O(n8529));
  invx  g07679(.a(n8421), .O(n8530));
  invx  g07680(.a(n8410), .O(n8531));
  andx  g07681(.a(n8423), .b(n8531), .O(n8532));
  orx   g07682(.a(n8532), .b(n8530), .O(n8533));
  andx  g07683(.a(n8532), .b(n8530), .O(n8534));
  invx  g07684(.a(n8534), .O(n8535));
  andx  g07685(.a(n8535), .b(n8533), .O(n8536));
  invx  g07686(.a(n8536), .O(n8537));
  andx  g07687(.a(n7931), .b(n3210), .O(n8538));
  invx  g07688(.a(n8404), .O(n8539));
  andx  g07689(.a(n8539), .b(n8403), .O(n8540));
  invx  g07690(.a(n8403), .O(n8541));
  andx  g07691(.a(n8404), .b(n8541), .O(n8542));
  orx   g07692(.a(n8542), .b(n8540), .O(n8543));
  andx  g07693(.a(n8543), .b(n8538), .O(n8544));
  andx  g07694(.a(n7791), .b(n3284), .O(n8545));
  andx  g07695(.a(n7938), .b(n3210), .O(n8546));
  andx  g07696(.a(n8546), .b(n8545), .O(n8547));
  andx  g07697(.a(n8547), .b(n8538), .O(n8548));
  andx  g07698(.a(n8547), .b(n8543), .O(n8549));
  orx   g07699(.a(n8549), .b(n8548), .O(n8550));
  orx   g07700(.a(n8550), .b(n8544), .O(n8551));
  andx  g07701(.a(n8551), .b(n7924), .O(n8552));
  invx  g07702(.a(n8405), .O(n8553));
  andx  g07703(.a(n8553), .b(n8396), .O(n8554));
  invx  g07704(.a(n8554), .O(n8555));
  orx   g07705(.a(n8553), .b(n8396), .O(n8556));
  andx  g07706(.a(n8556), .b(n8555), .O(n8557));
  andx  g07707(.a(n8397), .b(n8399), .O(n8558));
  orx   g07708(.a(n8558), .b(n8157), .O(n8559));
  andx  g07709(.a(n8559), .b(n8557), .O(n8560));
  invx  g07710(.a(n8560), .O(n8561));
  orx   g07711(.a(n8559), .b(n8557), .O(n8562));
  andx  g07712(.a(n8562), .b(n8561), .O(n8563));
  andx  g07713(.a(n7924), .b(n3210), .O(n8564));
  orx   g07714(.a(n8564), .b(n8551), .O(n8565));
  andx  g07715(.a(n8565), .b(n8563), .O(n8566));
  orx   g07716(.a(n8566), .b(n8552), .O(n8567));
  andx  g07717(.a(n8567), .b(n8537), .O(n8568));
  andx  g07718(.a(n7982), .b(n3210), .O(n8569));
  invx  g07719(.a(n8569), .O(n8570));
  invx  g07720(.a(n8567), .O(n8571));
  andx  g07721(.a(n8571), .b(n8536), .O(n8572));
  orx   g07722(.a(n8572), .b(n8570), .O(n8573));
  invx  g07723(.a(n8573), .O(n8574));
  orx   g07724(.a(n8574), .b(n8568), .O(n8575));
  andx  g07725(.a(n8575), .b(n8529), .O(n8576));
  orx   g07726(.a(n8575), .b(n8529), .O(n8577));
  andx  g07727(.a(n8062), .b(n3210), .O(n8578));
  andx  g07728(.a(n8578), .b(n8577), .O(n8579));
  orx   g07729(.a(n8579), .b(n8576), .O(n8580));
  andx  g07730(.a(n8580), .b(n8522), .O(n8581));
  andx  g07731(.a(n8131), .b(n3210), .O(n8582));
  orx   g07732(.a(n8580), .b(n8522), .O(n8583));
  andx  g07733(.a(n8583), .b(n8582), .O(n8584));
  orx   g07734(.a(n8584), .b(n8581), .O(n8585));
  andx  g07735(.a(n8585), .b(n8513), .O(n8586));
  orx   g07736(.a(n8585), .b(n8513), .O(n8587));
  andx  g07737(.a(n8220), .b(n3210), .O(n8588));
  andx  g07738(.a(n8588), .b(n8587), .O(n8589));
  orx   g07739(.a(n8589), .b(n8586), .O(n8590));
  andx  g07740(.a(n8590), .b(n8498), .O(n8591));
  andx  g07741(.a(n8351), .b(n3210), .O(n8592));
  orx   g07742(.a(n8590), .b(n8498), .O(n8593));
  andx  g07743(.a(n8593), .b(n8592), .O(n8594));
  orx   g07744(.a(n8594), .b(n8591), .O(n8595));
  andx  g07745(.a(n8595), .b(n8489), .O(n8596));
  orx   g07746(.a(n8595), .b(n8489), .O(n8597));
  andx  g07747(.a(n7864), .b(n8349), .O(n8598));
  andx  g07748(.a(n7858), .b(n7862), .O(n8599));
  andx  g07749(.a(n7859), .b(n7856), .O(n8600));
  orx   g07750(.a(n8600), .b(n8599), .O(n8601));
  andx  g07751(.a(n8601), .b(n7850), .O(n8602));
  orx   g07752(.a(n8602), .b(n8598), .O(n8603));
  andx  g07753(.a(n8603), .b(n3210), .O(n8604));
  andx  g07754(.a(n8604), .b(n8597), .O(n8605));
  orx   g07755(.a(n8605), .b(n8596), .O(n8606));
  andx  g07756(.a(n8606), .b(n7909), .O(n8607));
  invx  g07757(.a(n8596), .O(n8608));
  orx   g07758(.a(n8487), .b(n8484), .O(n8609));
  orx   g07759(.a(n8480), .b(n8345), .O(n8610));
  andx  g07760(.a(n8610), .b(n8609), .O(n8611));
  invx  g07761(.a(n8591), .O(n8612));
  invx  g07762(.a(n8592), .O(n8613));
  andx  g07763(.a(n8496), .b(n8370), .O(n8614));
  andx  g07764(.a(n8492), .b(n8449), .O(n8615));
  orx   g07765(.a(n8615), .b(n8614), .O(n8616));
  invx  g07766(.a(n8586), .O(n8617));
  orx   g07767(.a(n8511), .b(n8379), .O(n8618));
  orx   g07768(.a(n8507), .b(n8453), .O(n8619));
  andx  g07769(.a(n8619), .b(n8618), .O(n8620));
  invx  g07770(.a(n8581), .O(n8621));
  invx  g07771(.a(n8582), .O(n8622));
  orx   g07772(.a(n8520), .b(n8390), .O(n8623));
  orx   g07773(.a(n8516), .b(n8457), .O(n8624));
  andx  g07774(.a(n8624), .b(n8623), .O(n8625));
  invx  g07775(.a(n8576), .O(n8626));
  invx  g07776(.a(n8528), .O(n8627));
  orx   g07777(.a(n8627), .b(n8526), .O(n8628));
  invx  g07778(.a(n8568), .O(n8629));
  andx  g07779(.a(n8573), .b(n8629), .O(n8630));
  andx  g07780(.a(n8630), .b(n8628), .O(n8631));
  invx  g07781(.a(n8578), .O(n8632));
  orx   g07782(.a(n8632), .b(n8631), .O(n8633));
  andx  g07783(.a(n8633), .b(n8626), .O(n8634));
  andx  g07784(.a(n8634), .b(n8625), .O(n8635));
  orx   g07785(.a(n8635), .b(n8622), .O(n8636));
  andx  g07786(.a(n8636), .b(n8621), .O(n8637));
  andx  g07787(.a(n8637), .b(n8620), .O(n8638));
  invx  g07788(.a(n8588), .O(n8639));
  orx   g07789(.a(n8639), .b(n8638), .O(n8640));
  andx  g07790(.a(n8640), .b(n8617), .O(n8641));
  andx  g07791(.a(n8641), .b(n8616), .O(n8642));
  orx   g07792(.a(n8642), .b(n8613), .O(n8643));
  andx  g07793(.a(n8643), .b(n8612), .O(n8644));
  andx  g07794(.a(n8644), .b(n8611), .O(n8645));
  invx  g07795(.a(n8604), .O(n8646));
  orx   g07796(.a(n8646), .b(n8645), .O(n8647));
  andx  g07797(.a(n8647), .b(n8608), .O(n8648));
  andx  g07798(.a(n8648), .b(n7908), .O(n8649));
  orx   g07799(.a(n8649), .b(n8607), .O(n8650));
  andx  g07800(.a(n8220), .b(n3429), .O(n8651));
  orx   g07801(.a(n8294), .b(n8292), .O(n8652));
  orx   g07802(.a(n8288), .b(n8247), .O(n8653));
  andx  g07803(.a(n8653), .b(n8652), .O(n8654));
  andx  g07804(.a(n8304), .b(n8306), .O(n8655));
  andx  g07805(.a(n8310), .b(n8300), .O(n8656));
  orx   g07806(.a(n8656), .b(n8655), .O(n8657));
  andx  g07807(.a(n8657), .b(n8654), .O(n8658));
  orx   g07808(.a(n8313), .b(n8658), .O(n8663));
  andx  g07809(.a(n8663), .b(n8317), .O(n8664));
  invx  g07810(.a(n8664), .O(n8665));
  orx   g07811(.a(n8657), .b(n8654), .O(n8667));
  andx  g07812(.a(n8667), .b(n8315), .O(n8668));
  orx   g07813(.a(n8668), .b(n8327), .O(n8669));
  orx   g07814(.a(n8327), .b(n8318), .O(n8670));
  andx  g07815(.a(n8670), .b(n8669), .O(n8671));
  andx  g07816(.a(n8671), .b(n8665), .O(n8672));
  orx   g07817(.a(n8672), .b(n8651), .O(n8673));
  andx  g07818(.a(n8217), .b(n8211), .O(n8674));
  orx   g07819(.a(n8674), .b(n7849), .O(n8675));
  orx   g07820(.a(n8675), .b(n3297), .O(n8676));
  andx  g07821(.a(n8663), .b(n8322), .O(n8677));
  andx  g07822(.a(n8322), .b(n8317), .O(n8678));
  orx   g07823(.a(n8678), .b(n8677), .O(n8679));
  orx   g07824(.a(n8679), .b(n8664), .O(n8680));
  orx   g07825(.a(n8680), .b(n8676), .O(n8681));
  andx  g07826(.a(n8681), .b(n8673), .O(n8682));
  andx  g07827(.a(n7982), .b(n3645), .O(n8683));
  invx  g07828(.a(n8260), .O(n8684));
  orx   g07829(.a(n8282), .b(n8279), .O(n8685));
  orx   g07830(.a(n8275), .b(n8268), .O(n8686));
  andx  g07831(.a(n8686), .b(n8685), .O(n8687));
  orx   g07832(.a(n8687), .b(n8255), .O(n8688));
  andx  g07833(.a(n8688), .b(n8684), .O(n8689));
  andx  g07834(.a(n8689), .b(n8683), .O(n8690));
  orx   g07835(.a(n7916), .b(n4509), .O(n8691));
  andx  g07836(.a(n7924), .b(n3645), .O(n8692));
  orx   g07837(.a(n8692), .b(n8259), .O(n8693));
  andx  g07838(.a(n8284), .b(n8693), .O(n8694));
  orx   g07839(.a(n8694), .b(n8260), .O(n8695));
  andx  g07840(.a(n8695), .b(n8691), .O(n8696));
  orx   g07841(.a(n8696), .b(n8690), .O(n8697));
  andx  g07842(.a(n8266), .b(n8262), .O(n8698));
  invx  g07843(.a(n8698), .O(n8699));
  orx   g07844(.a(n8282), .b(n8263), .O(n8700));
  orx   g07845(.a(n8282), .b(n8265), .O(n8701));
  andx  g07846(.a(n8701), .b(n8700), .O(n8702));
  andx  g07847(.a(n8702), .b(n8699), .O(n8703));
  orx   g07848(.a(n8009), .b(n6829), .O(n8704));
  andx  g07849(.a(n8704), .b(n8703), .O(n8705));
  andx  g07850(.a(n8275), .b(n8266), .O(n8706));
  andx  g07851(.a(n8275), .b(n8262), .O(n8707));
  orx   g07852(.a(n8707), .b(n8706), .O(n8708));
  orx   g07853(.a(n8708), .b(n8698), .O(n8709));
  andx  g07854(.a(n8709), .b(n7924), .O(n8710));
  orx   g07855(.a(n8710), .b(n8705), .O(n8711));
  andx  g07856(.a(n8273), .b(n8269), .O(n8712));
  orx   g07857(.a(n7959), .b(n4062), .O(n8713));
  orx   g07858(.a(n8713), .b(n8712), .O(n8714));
  invx  g07859(.a(n8712), .O(n8715));
  andx  g07860(.a(n7931), .b(n4063), .O(n8716));
  orx   g07861(.a(n8716), .b(n8715), .O(n8717));
  andx  g07862(.a(n8717), .b(n8714), .O(n8718));
  andx  g07863(.a(n7791), .b(n4490), .O(n8719));
  andx  g07864(.a(n7938), .b(n4114), .O(n8720));
  orx   g07865(.a(n8720), .b(n8719), .O(n8721));
  andx  g07866(.a(n8720), .b(n8719), .O(n8722));
  invx  g07867(.a(n8722), .O(n8723));
  andx  g07868(.a(n8723), .b(n8721), .O(n8724));
  andx  g07869(.a(n8724), .b(n8718), .O(n8725));
  andx  g07870(.a(n8716), .b(n8715), .O(n8726));
  andx  g07871(.a(n8713), .b(n8712), .O(n8727));
  orx   g07872(.a(n8727), .b(n8726), .O(n8728));
  invx  g07873(.a(n8721), .O(n8729));
  orx   g07874(.a(n8722), .b(n8729), .O(n8730));
  andx  g07875(.a(n8730), .b(n8728), .O(n8731));
  orx   g07876(.a(n8731), .b(n8725), .O(n8732));
  andx  g07877(.a(n8732), .b(n8711), .O(n8733));
  orx   g07878(.a(n8732), .b(n8711), .O(n8734));
  invx  g07879(.a(n8734), .O(n8735));
  orx   g07880(.a(n8735), .b(n8733), .O(n8736));
  andx  g07881(.a(n8736), .b(n8697), .O(n8737));
  orx   g07882(.a(n8695), .b(n8691), .O(n8738));
  orx   g07883(.a(n8689), .b(n8683), .O(n8739));
  andx  g07884(.a(n8739), .b(n8738), .O(n8740));
  invx  g07885(.a(n8733), .O(n8741));
  andx  g07886(.a(n8734), .b(n8741), .O(n8742));
  andx  g07887(.a(n8742), .b(n8740), .O(n8743));
  orx   g07888(.a(n8743), .b(n8737), .O(n8744));
  orx   g07889(.a(n8299), .b(n4989), .O(n8745));
  andx  g07890(.a(n8245), .b(n8233), .O(n8746));
  orx   g07891(.a(n8245), .b(n8233), .O(n8747));
  andx  g07892(.a(n8747), .b(n8288), .O(n8748));
  orx   g07893(.a(n8748), .b(n8746), .O(n8749));
  andx  g07894(.a(n8749), .b(n8745), .O(n8750));
  andx  g07895(.a(n8062), .b(n3413), .O(n8751));
  invx  g07896(.a(n8746), .O(n8752));
  andx  g07897(.a(n8239), .b(n8241), .O(n8753));
  orx   g07898(.a(n8753), .b(n8294), .O(n8754));
  andx  g07899(.a(n8754), .b(n8752), .O(n8755));
  andx  g07900(.a(n8755), .b(n8751), .O(n8756));
  orx   g07901(.a(n8756), .b(n8750), .O(n8757));
  andx  g07902(.a(n8757), .b(n8744), .O(n8758));
  orx   g07903(.a(n8757), .b(n8744), .O(n8759));
  andx  g07904(.a(n8131), .b(n3171), .O(n8762));
  orx   g07905(.a(n8310), .b(n8296), .O(n8763));
  andx  g07906(.a(n8310), .b(n8296), .O(n8764));
  orx   g07907(.a(n8764), .b(n8300), .O(n8765));
  andx  g07908(.a(n8765), .b(n8763), .O(n8766));
  orx   g07909(.a(n8766), .b(n8762), .O(n8767));
  orx   g07910(.a(n8129), .b(n7835), .O(n8768));
  orx   g07911(.a(n7841), .b(n8124), .O(n8769));
  andx  g07912(.a(n8769), .b(n8768), .O(n8770));
  orx   g07913(.a(n8770), .b(n3418), .O(n8771));
  andx  g07914(.a(n8304), .b(n8654), .O(n8772));
  orx   g07915(.a(n8304), .b(n8654), .O(n8773));
  andx  g07916(.a(n8773), .b(n8306), .O(n8774));
  orx   g07917(.a(n8774), .b(n8772), .O(n8775));
  orx   g07918(.a(n8775), .b(n8771), .O(n8776));
  andx  g07919(.a(n8776), .b(n8767), .O(n8777));
  orx   g07920(.a(n8777), .b(n9700), .O(n8778));
  andx  g07921(.a(n8775), .b(n8771), .O(n8781));
  andx  g07922(.a(n8766), .b(n8762), .O(n8782));
  orx   g07923(.a(n8782), .b(n8781), .O(n8783));
  orx   g07924(.a(n8783), .b(n9711), .O(n8784));
  andx  g07925(.a(n8784), .b(n8778), .O(n8785));
  orx   g07926(.a(n8785), .b(n8682), .O(n8786));
  andx  g07927(.a(n8680), .b(n8676), .O(n8787));
  andx  g07928(.a(n8672), .b(n8651), .O(n8788));
  orx   g07929(.a(n8788), .b(n8787), .O(n8789));
  andx  g07930(.a(n8783), .b(n9711), .O(n8790));
  andx  g07931(.a(n8777), .b(n9700), .O(n8791));
  orx   g07932(.a(n8791), .b(n8790), .O(n8792));
  orx   g07933(.a(n8792), .b(n8789), .O(n8793));
  andx  g07934(.a(n8793), .b(n8786), .O(n8794));
  andx  g07935(.a(n8351), .b(n3180), .O(n8795));
  andx  g07936(.a(n8336), .b(n8229), .O(n8796));
  invx  g07937(.a(n8796), .O(n8797));
  andx  g07938(.a(n8343), .b(n8210), .O(n8798));
  orx   g07939(.a(n8798), .b(n8230), .O(n8799));
  andx  g07940(.a(n8799), .b(n8797), .O(n8800));
  orx   g07941(.a(n8800), .b(n8795), .O(n8801));
  invx  g07942(.a(n8795), .O(n8802));
  orx   g07943(.a(n8336), .b(n8229), .O(n8803));
  andx  g07944(.a(n8803), .b(n8221), .O(n8804));
  orx   g07945(.a(n8804), .b(n8796), .O(n8805));
  orx   g07946(.a(n8805), .b(n8802), .O(n8806));
  andx  g07947(.a(n8806), .b(n8801), .O(n8807));
  orx   g07948(.a(n8807), .b(n8794), .O(n8808));
  andx  g07949(.a(n8792), .b(n8789), .O(n8809));
  andx  g07950(.a(n8785), .b(n8682), .O(n8810));
  orx   g07951(.a(n8810), .b(n8809), .O(n8811));
  andx  g07952(.a(n8805), .b(n8802), .O(n8812));
  andx  g07953(.a(n8800), .b(n8795), .O(n8813));
  orx   g07954(.a(n8813), .b(n8812), .O(n8814));
  orx   g07955(.a(n8814), .b(n8811), .O(n8815));
  andx  g07956(.a(n8815), .b(n8808), .O(n8816));
  andx  g07957(.a(n8603), .b(n3284), .O(n8817));
  invx  g07958(.a(n8817), .O(n8818));
  andx  g07959(.a(n8352), .b(n8484), .O(n8819));
  andx  g07960(.a(n8444), .b(n8484), .O(n8820));
  andx  g07961(.a(n8444), .b(n8352), .O(n8821));
  orx   g07962(.a(n8821), .b(n8820), .O(n8822));
  orx   g07963(.a(n8822), .b(n8819), .O(n8823));
  andx  g07964(.a(n8823), .b(n8818), .O(n8824));
  invx  g07965(.a(n8819), .O(n8825));
  orx   g07966(.a(n8478), .b(n8345), .O(n8826));
  orx   g07967(.a(n8478), .b(n8353), .O(n8827));
  andx  g07968(.a(n8827), .b(n8826), .O(n8828));
  andx  g07969(.a(n8828), .b(n8825), .O(n8829));
  andx  g07970(.a(n8829), .b(n8817), .O(n8830));
  orx   g07971(.a(n8830), .b(n8824), .O(n8831));
  andx  g07972(.a(n9918), .b(n8650), .O(n8836));
  orx   g07973(.a(n8648), .b(n7908), .O(n8837));
  orx   g07974(.a(n8606), .b(n7909), .O(n8838));
  andx  g07975(.a(n8838), .b(n8837), .O(n8839));
  andx  g07976(.a(n9908), .b(n8839), .O(n8841));
  orx   g07977(.a(n8841), .b(n8836), .O(n8842));
  invx  g07978(.a(n7873), .O(n8843));
  andx  g07979(.a(n7738), .b(n5397), .O(n8844));
  andx  g07980(.a(n8844), .b(n7869), .O(n8845));
  andx  g07981(.a(n5777), .b(n7737), .O(n8846));
  andx  g07982(.a(n7868), .b(n7737), .O(n8847));
  orx   g07983(.a(n8847), .b(n8846), .O(n8848));
  orx   g07984(.a(n8848), .b(n8845), .O(n8849));
  orx   g07985(.a(n8849), .b(n8843), .O(n8850));
  orx   g07986(.a(n7879), .b(n7873), .O(n8851));
  andx  g07987(.a(n8851), .b(n8850), .O(n8852));
  andx  g07988(.a(n8852), .b(n3221), .O(n8853));
  andx  g07989(.a(n7907), .b(n3221), .O(n8854));
  orx   g07990(.a(n8646), .b(n8595), .O(n8855));
  orx   g07991(.a(n8604), .b(n8644), .O(n8856));
  andx  g07992(.a(n8856), .b(n8855), .O(n8857));
  andx  g07993(.a(n8857), .b(n8489), .O(n8858));
  andx  g07994(.a(n8604), .b(n8644), .O(n8859));
  andx  g07995(.a(n8646), .b(n8595), .O(n8860));
  orx   g07996(.a(n8860), .b(n8859), .O(n8861));
  andx  g07997(.a(n8861), .b(n8611), .O(n8862));
  orx   g07998(.a(n8862), .b(n8858), .O(n8863));
  andx  g07999(.a(n8863), .b(n8854), .O(n8864));
  invx  g08000(.a(n8864), .O(n8865));
  invx  g08001(.a(n8854), .O(n8866));
  andx  g08002(.a(n8613), .b(n8590), .O(n8867));
  andx  g08003(.a(n8592), .b(n8641), .O(n8868));
  orx   g08004(.a(n8868), .b(n8867), .O(n8869));
  andx  g08005(.a(n8869), .b(n8616), .O(n8870));
  orx   g08006(.a(n8592), .b(n8641), .O(n8871));
  orx   g08007(.a(n8613), .b(n8590), .O(n8872));
  andx  g08008(.a(n8872), .b(n8871), .O(n8873));
  andx  g08009(.a(n8873), .b(n8498), .O(n8874));
  orx   g08010(.a(n8874), .b(n8870), .O(n8875));
  andx  g08011(.a(n8639), .b(n8585), .O(n8876));
  andx  g08012(.a(n8588), .b(n8637), .O(n8877));
  orx   g08013(.a(n8877), .b(n8876), .O(n8878));
  andx  g08014(.a(n8878), .b(n8620), .O(n8879));
  orx   g08015(.a(n8588), .b(n8637), .O(n8880));
  orx   g08016(.a(n8639), .b(n8585), .O(n8881));
  andx  g08017(.a(n8881), .b(n8880), .O(n8882));
  andx  g08018(.a(n8882), .b(n8513), .O(n8883));
  orx   g08019(.a(n8883), .b(n8879), .O(n8884));
  orx   g08020(.a(n8582), .b(n8634), .O(n8885));
  orx   g08021(.a(n8622), .b(n8580), .O(n8886));
  andx  g08022(.a(n8886), .b(n8885), .O(n8887));
  orx   g08023(.a(n8887), .b(n8625), .O(n8888));
  andx  g08024(.a(n8622), .b(n8580), .O(n8889));
  andx  g08025(.a(n8582), .b(n8634), .O(n8890));
  orx   g08026(.a(n8890), .b(n8889), .O(n8891));
  orx   g08027(.a(n8891), .b(n8522), .O(n8892));
  andx  g08028(.a(n8892), .b(n8888), .O(n8893));
  andx  g08029(.a(n8632), .b(n8575), .O(n8894));
  andx  g08030(.a(n8578), .b(n8630), .O(n8895));
  orx   g08031(.a(n8895), .b(n8894), .O(n8896));
  andx  g08032(.a(n8896), .b(n8628), .O(n8897));
  orx   g08033(.a(n8578), .b(n8630), .O(n8898));
  orx   g08034(.a(n8632), .b(n8575), .O(n8899));
  andx  g08035(.a(n8899), .b(n8898), .O(n8900));
  andx  g08036(.a(n8900), .b(n8529), .O(n8901));
  orx   g08037(.a(n8901), .b(n8897), .O(n8902));
  andx  g08038(.a(n8570), .b(n8567), .O(n8903));
  andx  g08039(.a(n8569), .b(n8571), .O(n8904));
  orx   g08040(.a(n8904), .b(n8903), .O(n8905));
  andx  g08041(.a(n8905), .b(n8537), .O(n8906));
  invx  g08042(.a(n8906), .O(n8907));
  orx   g08043(.a(n8905), .b(n8537), .O(n8908));
  andx  g08044(.a(n8908), .b(n8907), .O(n8909));
  invx  g08045(.a(n8552), .O(n8910));
  andx  g08046(.a(n8565), .b(n8910), .O(n8911));
  invx  g08047(.a(n8911), .O(n8912));
  andx  g08048(.a(n8912), .b(n8563), .O(n8913));
  invx  g08049(.a(n8913), .O(n8914));
  orx   g08050(.a(n8912), .b(n8563), .O(n8915));
  andx  g08051(.a(n8915), .b(n8914), .O(n8916));
  invx  g08052(.a(n8916), .O(n8917));
  andx  g08053(.a(n7931), .b(n3221), .O(n8918));
  invx  g08054(.a(n8546), .O(n8919));
  andx  g08055(.a(n8919), .b(n8545), .O(n8920));
  invx  g08056(.a(n8545), .O(n8921));
  andx  g08057(.a(n8546), .b(n8921), .O(n8922));
  orx   g08058(.a(n8922), .b(n8920), .O(n8923));
  andx  g08059(.a(n8923), .b(n8918), .O(n8924));
  andx  g08060(.a(n7791), .b(n3210), .O(n8925));
  andx  g08061(.a(n7938), .b(n3221), .O(n8926));
  andx  g08062(.a(n8926), .b(n8925), .O(n8927));
  andx  g08063(.a(n8927), .b(n8918), .O(n8928));
  andx  g08064(.a(n8927), .b(n8923), .O(n8929));
  orx   g08065(.a(n8929), .b(n8928), .O(n8930));
  orx   g08066(.a(n8930), .b(n8924), .O(n8931));
  andx  g08067(.a(n8931), .b(n7924), .O(n8932));
  invx  g08068(.a(n8547), .O(n8933));
  andx  g08069(.a(n8933), .b(n8538), .O(n8934));
  invx  g08070(.a(n8934), .O(n8935));
  orx   g08071(.a(n8933), .b(n8538), .O(n8936));
  andx  g08072(.a(n8936), .b(n8935), .O(n8937));
  andx  g08073(.a(n8539), .b(n8541), .O(n8938));
  orx   g08074(.a(n8938), .b(n8405), .O(n8939));
  andx  g08075(.a(n8939), .b(n8937), .O(n8940));
  invx  g08076(.a(n8940), .O(n8941));
  orx   g08077(.a(n8939), .b(n8937), .O(n8942));
  andx  g08078(.a(n8942), .b(n8941), .O(n8943));
  andx  g08079(.a(n7924), .b(n3221), .O(n8944));
  orx   g08080(.a(n8944), .b(n8931), .O(n8945));
  andx  g08081(.a(n8945), .b(n8943), .O(n8946));
  orx   g08082(.a(n8946), .b(n8932), .O(n8947));
  andx  g08083(.a(n8947), .b(n8917), .O(n8948));
  andx  g08084(.a(n7982), .b(n3221), .O(n8949));
  invx  g08085(.a(n8949), .O(n8950));
  invx  g08086(.a(n8947), .O(n8951));
  andx  g08087(.a(n8951), .b(n8916), .O(n8952));
  orx   g08088(.a(n8952), .b(n8950), .O(n8953));
  invx  g08089(.a(n8953), .O(n8954));
  orx   g08090(.a(n8954), .b(n8948), .O(n8955));
  andx  g08091(.a(n8955), .b(n8909), .O(n8956));
  orx   g08092(.a(n8955), .b(n8909), .O(n8957));
  andx  g08093(.a(n8062), .b(n3221), .O(n8958));
  andx  g08094(.a(n8958), .b(n8957), .O(n8959));
  orx   g08095(.a(n8959), .b(n8956), .O(n8960));
  andx  g08096(.a(n8960), .b(n8902), .O(n8961));
  andx  g08097(.a(n8131), .b(n3221), .O(n8962));
  orx   g08098(.a(n8960), .b(n8902), .O(n8963));
  andx  g08099(.a(n8963), .b(n8962), .O(n8964));
  orx   g08100(.a(n8964), .b(n8961), .O(n8965));
  andx  g08101(.a(n8965), .b(n8893), .O(n8966));
  orx   g08102(.a(n8965), .b(n8893), .O(n8967));
  andx  g08103(.a(n8220), .b(n3221), .O(n8968));
  andx  g08104(.a(n8968), .b(n8967), .O(n8969));
  orx   g08105(.a(n8969), .b(n8966), .O(n8970));
  andx  g08106(.a(n8970), .b(n8884), .O(n8971));
  andx  g08107(.a(n8351), .b(n3221), .O(n8972));
  orx   g08108(.a(n8970), .b(n8884), .O(n8973));
  andx  g08109(.a(n8973), .b(n8972), .O(n8974));
  orx   g08110(.a(n8974), .b(n8971), .O(n8975));
  andx  g08111(.a(n8975), .b(n8875), .O(n8976));
  invx  g08112(.a(n8976), .O(n8977));
  orx   g08113(.a(n8873), .b(n8498), .O(n8978));
  orx   g08114(.a(n8869), .b(n8616), .O(n8979));
  andx  g08115(.a(n8979), .b(n8978), .O(n8980));
  invx  g08116(.a(n8971), .O(n8981));
  invx  g08117(.a(n8972), .O(n8982));
  orx   g08118(.a(n8882), .b(n8513), .O(n8983));
  orx   g08119(.a(n8878), .b(n8620), .O(n8984));
  andx  g08120(.a(n8984), .b(n8983), .O(n8985));
  invx  g08121(.a(n8966), .O(n8986));
  andx  g08122(.a(n8891), .b(n8522), .O(n8987));
  andx  g08123(.a(n8887), .b(n8625), .O(n8988));
  orx   g08124(.a(n8988), .b(n8987), .O(n8989));
  invx  g08125(.a(n8961), .O(n8990));
  invx  g08126(.a(n8962), .O(n8991));
  orx   g08127(.a(n8900), .b(n8529), .O(n8992));
  orx   g08128(.a(n8896), .b(n8628), .O(n8993));
  andx  g08129(.a(n8993), .b(n8992), .O(n8994));
  invx  g08130(.a(n8956), .O(n8995));
  invx  g08131(.a(n8909), .O(n8996));
  invx  g08132(.a(n8948), .O(n8997));
  andx  g08133(.a(n8953), .b(n8997), .O(n8998));
  andx  g08134(.a(n8998), .b(n8996), .O(n8999));
  invx  g08135(.a(n8958), .O(n9000));
  orx   g08136(.a(n9000), .b(n8999), .O(n9001));
  andx  g08137(.a(n9001), .b(n8995), .O(n9002));
  andx  g08138(.a(n9002), .b(n8994), .O(n9003));
  orx   g08139(.a(n9003), .b(n8991), .O(n9004));
  andx  g08140(.a(n9004), .b(n8990), .O(n9005));
  andx  g08141(.a(n9005), .b(n8989), .O(n9006));
  invx  g08142(.a(n8968), .O(n9007));
  orx   g08143(.a(n9007), .b(n9006), .O(n9008));
  andx  g08144(.a(n9008), .b(n8986), .O(n9009));
  andx  g08145(.a(n9009), .b(n8985), .O(n9010));
  orx   g08146(.a(n9010), .b(n8982), .O(n9011));
  andx  g08147(.a(n9011), .b(n8981), .O(n9012));
  andx  g08148(.a(n9012), .b(n8980), .O(n9013));
  andx  g08149(.a(n8603), .b(n3221), .O(n9014));
  invx  g08150(.a(n9014), .O(n9015));
  orx   g08151(.a(n9015), .b(n9013), .O(n9016));
  andx  g08152(.a(n9016), .b(n8977), .O(n9017));
  orx   g08153(.a(n9017), .b(n8866), .O(n9018));
  orx   g08154(.a(n8861), .b(n8611), .O(n9019));
  orx   g08155(.a(n8857), .b(n8489), .O(n9020));
  andx  g08156(.a(n9020), .b(n9019), .O(n9021));
  orx   g08157(.a(n9017), .b(n9021), .O(n9022));
  andx  g08158(.a(n9022), .b(n9018), .O(n9023));
  andx  g08159(.a(n9023), .b(n8865), .O(n9024));
  orx   g08160(.a(n9024), .b(n8853), .O(n9025));
  invx  g08161(.a(n8853), .O(n9026));
  orx   g08162(.a(n8975), .b(n8875), .O(n9027));
  andx  g08163(.a(n9014), .b(n9027), .O(n9028));
  orx   g08164(.a(n9028), .b(n8976), .O(n9029));
  andx  g08165(.a(n9029), .b(n8854), .O(n9030));
  andx  g08166(.a(n9029), .b(n8863), .O(n9031));
  orx   g08167(.a(n9031), .b(n9030), .O(n9032));
  orx   g08168(.a(n9032), .b(n8864), .O(n9033));
  orx   g08169(.a(n9033), .b(n9026), .O(n9034));
  andx  g08170(.a(n9034), .b(n9025), .O(n9035));
  orx   g08171(.a(n9035), .b(n8842), .O(n9036));
  orx   g08172(.a(n9908), .b(n8839), .O(n9037));
  orx   g08173(.a(n9918), .b(n8650), .O(n9038));
  andx  g08174(.a(n9038), .b(n9037), .O(n9039));
  andx  g08175(.a(n9033), .b(n9026), .O(n9040));
  andx  g08176(.a(n9024), .b(n8853), .O(n9041));
  orx   g08177(.a(n9041), .b(n9040), .O(n9042));
  orx   g08178(.a(n9042), .b(n9039), .O(n9043));
  andx  g08179(.a(n9043), .b(n9036), .O(n9044));
  orx   g08180(.a(n7761), .b(n7760), .O(n9045));
  orx   g08181(.a(n7757), .b(n7734), .O(n9046));
  andx  g08182(.a(n9046), .b(n9045), .O(n9047));
  orx   g08183(.a(n8850), .b(n9047), .O(n9048));
  orx   g08184(.a(n7880), .b(n7763), .O(n9049));
  andx  g08185(.a(n9049), .b(n9048), .O(n9050));
  andx  g08186(.a(n9050), .b(n3230), .O(n9051));
  invx  g08187(.a(n9051), .O(n9052));
  orx   g08188(.a(n9029), .b(n8854), .O(n9060));
  andx  g08189(.a(n9060), .b(n9018), .O(n9061));
  andx  g08190(.a(n9061), .b(n9021), .O(n9062));
  andx  g08191(.a(n9017), .b(n8866), .O(n9064));
  orx   g08192(.a(n9064), .b(n9030), .O(n9065));
  andx  g08193(.a(n9065), .b(n8863), .O(n9066));
  orx   g08194(.a(n9066), .b(n9062), .O(n9067));
  andx  g08195(.a(n9015), .b(n8975), .O(n9068));
  andx  g08196(.a(n9014), .b(n9012), .O(n9069));
  orx   g08197(.a(n9069), .b(n9068), .O(n9070));
  andx  g08198(.a(n9070), .b(n8980), .O(n9071));
  orx   g08199(.a(n9014), .b(n9012), .O(n9072));
  orx   g08200(.a(n9015), .b(n8975), .O(n9073));
  andx  g08201(.a(n9073), .b(n9072), .O(n9074));
  andx  g08202(.a(n9074), .b(n8875), .O(n9075));
  orx   g08203(.a(n9075), .b(n9071), .O(n9076));
  andx  g08204(.a(n8982), .b(n8970), .O(n9077));
  andx  g08205(.a(n8972), .b(n9009), .O(n9078));
  orx   g08206(.a(n9078), .b(n9077), .O(n9079));
  andx  g08207(.a(n9079), .b(n8985), .O(n9080));
  orx   g08208(.a(n8972), .b(n9009), .O(n9081));
  orx   g08209(.a(n8982), .b(n8970), .O(n9082));
  andx  g08210(.a(n9082), .b(n9081), .O(n9083));
  andx  g08211(.a(n9083), .b(n8884), .O(n9084));
  orx   g08212(.a(n9084), .b(n9080), .O(n9085));
  orx   g08213(.a(n9007), .b(n8965), .O(n9086));
  orx   g08214(.a(n8968), .b(n9005), .O(n9087));
  andx  g08215(.a(n9087), .b(n9086), .O(n9088));
  orx   g08216(.a(n9088), .b(n8989), .O(n9089));
  andx  g08217(.a(n8968), .b(n9005), .O(n9090));
  andx  g08218(.a(n9007), .b(n8965), .O(n9091));
  orx   g08219(.a(n9091), .b(n9090), .O(n9092));
  orx   g08220(.a(n9092), .b(n8893), .O(n9093));
  andx  g08221(.a(n9093), .b(n9089), .O(n9094));
  andx  g08222(.a(n8991), .b(n8960), .O(n9095));
  andx  g08223(.a(n8962), .b(n9002), .O(n9096));
  orx   g08224(.a(n9096), .b(n9095), .O(n9097));
  andx  g08225(.a(n9097), .b(n8994), .O(n9098));
  orx   g08226(.a(n8962), .b(n9002), .O(n9099));
  orx   g08227(.a(n8991), .b(n8960), .O(n9100));
  andx  g08228(.a(n9100), .b(n9099), .O(n9101));
  andx  g08229(.a(n9101), .b(n8902), .O(n9102));
  orx   g08230(.a(n9102), .b(n9098), .O(n9103));
  andx  g08231(.a(n9000), .b(n8955), .O(n9104));
  andx  g08232(.a(n8958), .b(n8998), .O(n9105));
  orx   g08233(.a(n9105), .b(n9104), .O(n9106));
  andx  g08234(.a(n9106), .b(n8996), .O(n9107));
  orx   g08235(.a(n8958), .b(n8998), .O(n9108));
  orx   g08236(.a(n9000), .b(n8955), .O(n9109));
  andx  g08237(.a(n9109), .b(n9108), .O(n9110));
  andx  g08238(.a(n9110), .b(n8909), .O(n9111));
  orx   g08239(.a(n9111), .b(n9107), .O(n9112));
  andx  g08240(.a(n8950), .b(n8947), .O(n9113));
  andx  g08241(.a(n8949), .b(n8951), .O(n9114));
  orx   g08242(.a(n9114), .b(n9113), .O(n9115));
  andx  g08243(.a(n9115), .b(n8917), .O(n9116));
  invx  g08244(.a(n9116), .O(n9117));
  orx   g08245(.a(n9115), .b(n8917), .O(n9118));
  andx  g08246(.a(n9118), .b(n9117), .O(n9119));
  invx  g08247(.a(n8932), .O(n9120));
  andx  g08248(.a(n8945), .b(n9120), .O(n9121));
  invx  g08249(.a(n9121), .O(n9122));
  andx  g08250(.a(n9122), .b(n8943), .O(n9123));
  invx  g08251(.a(n9123), .O(n9124));
  orx   g08252(.a(n9122), .b(n8943), .O(n9125));
  andx  g08253(.a(n9125), .b(n9124), .O(n9126));
  invx  g08254(.a(n9126), .O(n9127));
  andx  g08255(.a(n7931), .b(n3230), .O(n9128));
  invx  g08256(.a(n8926), .O(n9129));
  andx  g08257(.a(n9129), .b(n8925), .O(n9130));
  invx  g08258(.a(n8925), .O(n9131));
  andx  g08259(.a(n8926), .b(n9131), .O(n9132));
  orx   g08260(.a(n9132), .b(n9130), .O(n9133));
  andx  g08261(.a(n9133), .b(n9128), .O(n9134));
  andx  g08262(.a(n7791), .b(n3221), .O(n9135));
  andx  g08263(.a(n7938), .b(n3230), .O(n9136));
  andx  g08264(.a(n9136), .b(n9135), .O(n9137));
  andx  g08265(.a(n9137), .b(n9128), .O(n9138));
  andx  g08266(.a(n9137), .b(n9133), .O(n9139));
  orx   g08267(.a(n9139), .b(n9138), .O(n9140));
  orx   g08268(.a(n9140), .b(n9134), .O(n9141));
  andx  g08269(.a(n9141), .b(n7924), .O(n9142));
  invx  g08270(.a(n8927), .O(n9143));
  andx  g08271(.a(n9143), .b(n8918), .O(n9144));
  invx  g08272(.a(n9144), .O(n9145));
  orx   g08273(.a(n9143), .b(n8918), .O(n9146));
  andx  g08274(.a(n9146), .b(n9145), .O(n9147));
  andx  g08275(.a(n8919), .b(n8921), .O(n9148));
  orx   g08276(.a(n9148), .b(n8547), .O(n9149));
  andx  g08277(.a(n9149), .b(n9147), .O(n9150));
  invx  g08278(.a(n9150), .O(n9151));
  orx   g08279(.a(n9149), .b(n9147), .O(n9152));
  andx  g08280(.a(n9152), .b(n9151), .O(n9153));
  andx  g08281(.a(n7924), .b(n3230), .O(n9154));
  orx   g08282(.a(n9154), .b(n9141), .O(n9155));
  andx  g08283(.a(n9155), .b(n9153), .O(n9156));
  orx   g08284(.a(n9156), .b(n9142), .O(n9157));
  andx  g08285(.a(n9157), .b(n9127), .O(n9158));
  invx  g08286(.a(n9158), .O(n9159));
  andx  g08287(.a(n7982), .b(n3230), .O(n9160));
  invx  g08288(.a(n9160), .O(n9161));
  invx  g08289(.a(n9157), .O(n9162));
  andx  g08290(.a(n9162), .b(n9126), .O(n9163));
  orx   g08291(.a(n9163), .b(n9161), .O(n9164));
  andx  g08292(.a(n9164), .b(n9159), .O(n9165));
  invx  g08293(.a(n9165), .O(n9166));
  andx  g08294(.a(n9166), .b(n9119), .O(n9167));
  orx   g08295(.a(n9166), .b(n9119), .O(n9168));
  andx  g08296(.a(n8062), .b(n3230), .O(n9169));
  andx  g08297(.a(n9169), .b(n9168), .O(n9170));
  orx   g08298(.a(n9170), .b(n9167), .O(n9171));
  andx  g08299(.a(n9171), .b(n9112), .O(n9172));
  andx  g08300(.a(n8131), .b(n3230), .O(n9173));
  orx   g08301(.a(n9171), .b(n9112), .O(n9174));
  andx  g08302(.a(n9174), .b(n9173), .O(n9175));
  orx   g08303(.a(n9175), .b(n9172), .O(n9176));
  andx  g08304(.a(n9176), .b(n9103), .O(n9177));
  orx   g08305(.a(n9176), .b(n9103), .O(n9178));
  andx  g08306(.a(n8220), .b(n3230), .O(n9179));
  andx  g08307(.a(n9179), .b(n9178), .O(n9180));
  orx   g08308(.a(n9180), .b(n9177), .O(n9181));
  andx  g08309(.a(n9181), .b(n9094), .O(n9182));
  andx  g08310(.a(n8351), .b(n3230), .O(n9183));
  orx   g08311(.a(n9181), .b(n9094), .O(n9184));
  andx  g08312(.a(n9184), .b(n9183), .O(n9185));
  orx   g08313(.a(n9185), .b(n9182), .O(n9186));
  andx  g08314(.a(n9186), .b(n9085), .O(n9187));
  orx   g08315(.a(n9186), .b(n9085), .O(n9188));
  andx  g08316(.a(n8603), .b(n3230), .O(n9189));
  andx  g08317(.a(n9189), .b(n9188), .O(n9190));
  orx   g08318(.a(n9190), .b(n9187), .O(n9191));
  andx  g08319(.a(n9191), .b(n9076), .O(n9192));
  andx  g08320(.a(n7907), .b(n3230), .O(n9193));
  orx   g08321(.a(n9191), .b(n9076), .O(n9194));
  andx  g08322(.a(n9194), .b(n9193), .O(n9195));
  orx   g08323(.a(n9195), .b(n9192), .O(n9196));
  andx  g08324(.a(n9196), .b(n9067), .O(n9197));
  orx   g08325(.a(n9196), .b(n9067), .O(n9198));
  andx  g08326(.a(n8852), .b(n3230), .O(n9199));
  andx  g08327(.a(n9199), .b(n9198), .O(n9200));
  orx   g08328(.a(n9200), .b(n9197), .O(n9201));
  andx  g08329(.a(n9201), .b(n9052), .O(n9202));
  invx  g08330(.a(n9197), .O(n9203));
  orx   g08331(.a(n9065), .b(n8863), .O(n9204));
  orx   g08332(.a(n9061), .b(n9021), .O(n9205));
  andx  g08333(.a(n9205), .b(n9204), .O(n9206));
  invx  g08334(.a(n9192), .O(n9207));
  invx  g08335(.a(n9193), .O(n9208));
  orx   g08336(.a(n9074), .b(n8875), .O(n9209));
  orx   g08337(.a(n9070), .b(n8980), .O(n9210));
  andx  g08338(.a(n9210), .b(n9209), .O(n9211));
  invx  g08339(.a(n9187), .O(n9212));
  orx   g08340(.a(n9083), .b(n8884), .O(n9213));
  orx   g08341(.a(n9079), .b(n8985), .O(n9214));
  andx  g08342(.a(n9214), .b(n9213), .O(n9215));
  invx  g08343(.a(n9182), .O(n9216));
  invx  g08344(.a(n9183), .O(n9217));
  andx  g08345(.a(n9092), .b(n8893), .O(n9218));
  andx  g08346(.a(n9088), .b(n8989), .O(n9219));
  orx   g08347(.a(n9219), .b(n9218), .O(n9220));
  invx  g08348(.a(n9177), .O(n9221));
  orx   g08349(.a(n9101), .b(n8902), .O(n9222));
  orx   g08350(.a(n9097), .b(n8994), .O(n9223));
  andx  g08351(.a(n9223), .b(n9222), .O(n9224));
  invx  g08352(.a(n9172), .O(n9225));
  invx  g08353(.a(n9173), .O(n9226));
  orx   g08354(.a(n9110), .b(n8909), .O(n9227));
  orx   g08355(.a(n9106), .b(n8996), .O(n9228));
  andx  g08356(.a(n9228), .b(n9227), .O(n9229));
  invx  g08357(.a(n9167), .O(n9230));
  invx  g08358(.a(n9119), .O(n9231));
  andx  g08359(.a(n9165), .b(n9231), .O(n9232));
  invx  g08360(.a(n9169), .O(n9233));
  orx   g08361(.a(n9233), .b(n9232), .O(n9234));
  andx  g08362(.a(n9234), .b(n9230), .O(n9235));
  andx  g08363(.a(n9235), .b(n9229), .O(n9236));
  orx   g08364(.a(n9236), .b(n9226), .O(n9237));
  andx  g08365(.a(n9237), .b(n9225), .O(n9238));
  andx  g08366(.a(n9238), .b(n9224), .O(n9239));
  invx  g08367(.a(n9179), .O(n9240));
  orx   g08368(.a(n9240), .b(n9239), .O(n9241));
  andx  g08369(.a(n9241), .b(n9221), .O(n9242));
  andx  g08370(.a(n9242), .b(n9220), .O(n9243));
  orx   g08371(.a(n9243), .b(n9217), .O(n9244));
  andx  g08372(.a(n9244), .b(n9216), .O(n9245));
  andx  g08373(.a(n9245), .b(n9215), .O(n9246));
  invx  g08374(.a(n9189), .O(n9247));
  orx   g08375(.a(n9247), .b(n9246), .O(n9248));
  andx  g08376(.a(n9248), .b(n9212), .O(n9249));
  andx  g08377(.a(n9249), .b(n9211), .O(n9250));
  orx   g08378(.a(n9250), .b(n9208), .O(n9251));
  andx  g08379(.a(n9251), .b(n9207), .O(n9252));
  andx  g08380(.a(n9252), .b(n9206), .O(n9253));
  invx  g08381(.a(n9199), .O(n9254));
  orx   g08382(.a(n9254), .b(n9253), .O(n9255));
  andx  g08383(.a(n9255), .b(n9203), .O(n9256));
  andx  g08384(.a(n9256), .b(n9051), .O(n9257));
  orx   g08385(.a(n9257), .b(n9202), .O(n9258));
  andx  g08386(.a(n9258), .b(n9044), .O(n9259));
  invx  g08387(.a(n9259), .O(n9260));
  orx   g08388(.a(n9258), .b(n9044), .O(n9261));
  andx  g08389(.a(n9261), .b(n9260), .O(n9262));
  andx  g08390(.a(n7889), .b(n9048), .O(n9263));
  invx  g08391(.a(n9263), .O(n9264));
  orx   g08392(.a(n7889), .b(n9048), .O(n9265));
  andx  g08393(.a(n9265), .b(n9264), .O(n9266));
  invx  g08394(.a(n9266), .O(n9267));
  andx  g08395(.a(n9267), .b(n3258), .O(n9268));
  andx  g08396(.a(n9254), .b(n9196), .O(n9269));
  andx  g08397(.a(n9199), .b(n9252), .O(n9270));
  orx   g08398(.a(n9270), .b(n9269), .O(n9271));
  andx  g08399(.a(n9271), .b(n9206), .O(n9272));
  orx   g08400(.a(n9271), .b(n9206), .O(n9273));
  invx  g08401(.a(n9273), .O(n9274));
  orx   g08402(.a(n9274), .b(n9272), .O(n9275));
  andx  g08403(.a(n9208), .b(n9249), .O(n9276));
  andx  g08404(.a(n9193), .b(n9191), .O(n9277));
  orx   g08405(.a(n9277), .b(n9276), .O(n9278));
  orx   g08406(.a(n9278), .b(n9076), .O(n9279));
  invx  g08407(.a(n9279), .O(n9280));
  andx  g08408(.a(n9278), .b(n9076), .O(n9281));
  orx   g08409(.a(n9281), .b(n9280), .O(n9282));
  andx  g08410(.a(n9217), .b(n9181), .O(n9283));
  andx  g08411(.a(n9183), .b(n9242), .O(n9284));
  orx   g08412(.a(n9284), .b(n9283), .O(n9285));
  andx  g08413(.a(n9285), .b(n9220), .O(n9286));
  orx   g08414(.a(n9285), .b(n9220), .O(n9287));
  invx  g08415(.a(n9287), .O(n9288));
  orx   g08416(.a(n9288), .b(n9286), .O(n9289));
  andx  g08417(.a(n9226), .b(n9171), .O(n9290));
  andx  g08418(.a(n9173), .b(n9235), .O(n9291));
  orx   g08419(.a(n9291), .b(n9290), .O(n9292));
  andx  g08420(.a(n9292), .b(n9112), .O(n9293));
  invx  g08421(.a(n9293), .O(n9294));
  orx   g08422(.a(n9292), .b(n9112), .O(n9295));
  andx  g08423(.a(n9295), .b(n9294), .O(n9296));
  andx  g08424(.a(n9161), .b(n9157), .O(n9297));
  andx  g08425(.a(n9160), .b(n9162), .O(n9298));
  orx   g08426(.a(n9298), .b(n9297), .O(n9299));
  andx  g08427(.a(n9299), .b(n9127), .O(n9300));
  invx  g08428(.a(n9300), .O(n9301));
  orx   g08429(.a(n9299), .b(n9127), .O(n9302));
  andx  g08430(.a(n9302), .b(n9301), .O(n9303));
  invx  g08431(.a(n9142), .O(n9304));
  andx  g08432(.a(n9155), .b(n9304), .O(n9305));
  invx  g08433(.a(n9305), .O(n9306));
  andx  g08434(.a(n9306), .b(n9153), .O(n9307));
  invx  g08435(.a(n9307), .O(n9308));
  orx   g08436(.a(n9306), .b(n9153), .O(n9309));
  andx  g08437(.a(n9309), .b(n9308), .O(n9310));
  invx  g08438(.a(n9310), .O(n9311));
  invx  g08439(.a(n9137), .O(n9312));
  andx  g08440(.a(n9312), .b(n9128), .O(n9313));
  invx  g08441(.a(n9313), .O(n9314));
  orx   g08442(.a(n9312), .b(n9128), .O(n9315));
  andx  g08443(.a(n9315), .b(n9314), .O(n9316));
  andx  g08444(.a(n9129), .b(n9131), .O(n9317));
  orx   g08445(.a(n9317), .b(n8927), .O(n9318));
  andx  g08446(.a(n9318), .b(n9316), .O(n9319));
  invx  g08447(.a(n9319), .O(n9320));
  orx   g08448(.a(n9318), .b(n9316), .O(n9321));
  andx  g08449(.a(n9321), .b(n9320), .O(n9322));
  andx  g08450(.a(n7938), .b(n3258), .O(n9323));
  andx  g08451(.a(n9323), .b(n7791), .O(n9324));
  andx  g08452(.a(n9324), .b(n3230), .O(n9325));
  andx  g08453(.a(n9325), .b(n7931), .O(n9326));
  orx   g08454(.a(n9136), .b(n9135), .O(n9327));
  andx  g08455(.a(n9327), .b(n9312), .O(n9328));
  andx  g08456(.a(n7931), .b(n3258), .O(n9329));
  orx   g08457(.a(n9329), .b(n9325), .O(n9330));
  andx  g08458(.a(n9330), .b(n9328), .O(n9331));
  orx   g08459(.a(n9331), .b(n9326), .O(n9332));
  andx  g08460(.a(n9332), .b(n9322), .O(n9333));
  invx  g08461(.a(n9333), .O(n9334));
  invx  g08462(.a(n9322), .O(n9335));
  invx  g08463(.a(n9332), .O(n9336));
  andx  g08464(.a(n9336), .b(n9335), .O(n9337));
  andx  g08465(.a(n7924), .b(n3258), .O(n9338));
  invx  g08466(.a(n9338), .O(n9339));
  orx   g08467(.a(n9339), .b(n9337), .O(n9340));
  andx  g08468(.a(n9340), .b(n9334), .O(n9341));
  invx  g08469(.a(n9341), .O(n9342));
  andx  g08470(.a(n9342), .b(n9311), .O(n9343));
  invx  g08471(.a(n9343), .O(n9344));
  andx  g08472(.a(n9341), .b(n9310), .O(n9345));
  andx  g08473(.a(n7982), .b(n3258), .O(n9346));
  invx  g08474(.a(n9346), .O(n9347));
  orx   g08475(.a(n9347), .b(n9345), .O(n9348));
  andx  g08476(.a(n9348), .b(n9344), .O(n9349));
  invx  g08477(.a(n9349), .O(n9350));
  andx  g08478(.a(n9350), .b(n9303), .O(n9351));
  invx  g08479(.a(n9351), .O(n9352));
  invx  g08480(.a(n9303), .O(n9353));
  andx  g08481(.a(n9349), .b(n9353), .O(n9354));
  andx  g08482(.a(n8062), .b(n3258), .O(n9355));
  invx  g08483(.a(n9355), .O(n9356));
  orx   g08484(.a(n9356), .b(n9354), .O(n9357));
  andx  g08485(.a(n9357), .b(n9352), .O(n9358));
  invx  g08486(.a(n9358), .O(n9359));
  andx  g08487(.a(n9359), .b(n8131), .O(n9360));
  invx  g08488(.a(n9360), .O(n9361));
  andx  g08489(.a(n9233), .b(n9166), .O(n9362));
  andx  g08490(.a(n9169), .b(n9165), .O(n9363));
  orx   g08491(.a(n9363), .b(n9362), .O(n9364));
  andx  g08492(.a(n9364), .b(n9231), .O(n9365));
  invx  g08493(.a(n9365), .O(n9366));
  orx   g08494(.a(n9364), .b(n9231), .O(n9367));
  andx  g08495(.a(n9367), .b(n9366), .O(n9368));
  andx  g08496(.a(n8131), .b(n3258), .O(n9369));
  invx  g08497(.a(n9369), .O(n9370));
  andx  g08498(.a(n9370), .b(n9358), .O(n9371));
  orx   g08499(.a(n9371), .b(n9368), .O(n9372));
  andx  g08500(.a(n9372), .b(n9361), .O(n9373));
  invx  g08501(.a(n9373), .O(n9374));
  andx  g08502(.a(n9374), .b(n9296), .O(n9375));
  orx   g08503(.a(n9374), .b(n9296), .O(n9376));
  andx  g08504(.a(n8220), .b(n3258), .O(n9377));
  andx  g08505(.a(n9377), .b(n9376), .O(n9378));
  orx   g08506(.a(n9378), .b(n9375), .O(n9379));
  andx  g08507(.a(n9379), .b(n8351), .O(n9380));
  andx  g08508(.a(n9240), .b(n9176), .O(n9381));
  andx  g08509(.a(n9179), .b(n9238), .O(n9382));
  orx   g08510(.a(n9382), .b(n9381), .O(n9383));
  andx  g08511(.a(n9383), .b(n9224), .O(n9384));
  invx  g08512(.a(n9384), .O(n9385));
  orx   g08513(.a(n9383), .b(n9224), .O(n9386));
  andx  g08514(.a(n9386), .b(n9385), .O(n9387));
  invx  g08515(.a(n9387), .O(n9388));
  andx  g08516(.a(n8351), .b(n3258), .O(n9389));
  orx   g08517(.a(n9389), .b(n9379), .O(n9390));
  andx  g08518(.a(n9390), .b(n9388), .O(n9391));
  orx   g08519(.a(n9391), .b(n9380), .O(n9392));
  andx  g08520(.a(n9392), .b(n9289), .O(n9393));
  orx   g08521(.a(n9392), .b(n9289), .O(n9394));
  andx  g08522(.a(n8603), .b(n3258), .O(n9395));
  andx  g08523(.a(n9395), .b(n9394), .O(n9396));
  orx   g08524(.a(n9396), .b(n9393), .O(n9397));
  andx  g08525(.a(n9397), .b(n7907), .O(n9398));
  andx  g08526(.a(n9247), .b(n9245), .O(n9399));
  andx  g08527(.a(n9189), .b(n9186), .O(n9400));
  orx   g08528(.a(n9400), .b(n9399), .O(n9401));
  invx  g08529(.a(n9401), .O(n9402));
  andx  g08530(.a(n9402), .b(n9215), .O(n9403));
  andx  g08531(.a(n9401), .b(n9085), .O(n9404));
  orx   g08532(.a(n9404), .b(n9403), .O(n9405));
  andx  g08533(.a(n7907), .b(n3258), .O(n9406));
  orx   g08534(.a(n9406), .b(n9397), .O(n9407));
  andx  g08535(.a(n9407), .b(n9405), .O(n9408));
  orx   g08536(.a(n9408), .b(n9398), .O(n9409));
  andx  g08537(.a(n9409), .b(n9282), .O(n9410));
  orx   g08538(.a(n9409), .b(n9282), .O(n9411));
  andx  g08539(.a(n8852), .b(n3258), .O(n9412));
  andx  g08540(.a(n9412), .b(n9411), .O(n9413));
  orx   g08541(.a(n9413), .b(n9410), .O(n9414));
  andx  g08542(.a(n9414), .b(n9275), .O(n9415));
  orx   g08543(.a(n9414), .b(n9275), .O(n9416));
  andx  g08544(.a(n9050), .b(n3258), .O(n9417));
  andx  g08545(.a(n9417), .b(n9416), .O(n9418));
  orx   g08546(.a(n9418), .b(n9415), .O(n9419));
  andx  g08547(.a(n9419), .b(n9268), .O(n9420));
  invx  g08548(.a(n9268), .O(n9421));
  invx  g08549(.a(n9415), .O(n9422));
  invx  g08550(.a(n9272), .O(n9423));
  andx  g08551(.a(n9273), .b(n9423), .O(n9424));
  invx  g08552(.a(n9410), .O(n9425));
  invx  g08553(.a(n9281), .O(n9426));
  andx  g08554(.a(n9426), .b(n9279), .O(n9427));
  invx  g08555(.a(n9398), .O(n9428));
  invx  g08556(.a(n9405), .O(n9429));
  invx  g08557(.a(n9393), .O(n9430));
  invx  g08558(.a(n9286), .O(n9431));
  andx  g08559(.a(n9287), .b(n9431), .O(n9432));
  invx  g08560(.a(n9380), .O(n9433));
  invx  g08561(.a(n9375), .O(n9434));
  invx  g08562(.a(n9295), .O(n9435));
  orx   g08563(.a(n9435), .b(n9293), .O(n9436));
  andx  g08564(.a(n9373), .b(n9436), .O(n9437));
  invx  g08565(.a(n9377), .O(n9438));
  orx   g08566(.a(n9438), .b(n9437), .O(n9439));
  andx  g08567(.a(n9439), .b(n9434), .O(n9440));
  invx  g08568(.a(n9389), .O(n9441));
  andx  g08569(.a(n9441), .b(n9440), .O(n9442));
  orx   g08570(.a(n9442), .b(n9387), .O(n9443));
  andx  g08571(.a(n9443), .b(n9433), .O(n9444));
  andx  g08572(.a(n9444), .b(n9432), .O(n9445));
  invx  g08573(.a(n9395), .O(n9446));
  orx   g08574(.a(n9446), .b(n9445), .O(n9447));
  andx  g08575(.a(n9447), .b(n9430), .O(n9448));
  invx  g08576(.a(n9406), .O(n9449));
  andx  g08577(.a(n9449), .b(n9448), .O(n9450));
  orx   g08578(.a(n9450), .b(n9429), .O(n9451));
  andx  g08579(.a(n9451), .b(n9428), .O(n9452));
  andx  g08580(.a(n9452), .b(n9427), .O(n9453));
  invx  g08581(.a(n9412), .O(n9454));
  orx   g08582(.a(n9454), .b(n9453), .O(n9455));
  andx  g08583(.a(n9455), .b(n9425), .O(n9456));
  andx  g08584(.a(n9456), .b(n9424), .O(n9457));
  invx  g08585(.a(n9417), .O(n9458));
  orx   g08586(.a(n9458), .b(n9457), .O(n9459));
  andx  g08587(.a(n9459), .b(n9422), .O(n9460));
  andx  g08588(.a(n9460), .b(n9421), .O(n9461));
  orx   g08589(.a(n9461), .b(n9420), .O(n9462));
  andx  g08590(.a(n9462), .b(n9262), .O(n9463));
  invx  g08591(.a(n9463), .O(n9464));
  orx   g08592(.a(n9462), .b(n9262), .O(n9465));
  andx  g08593(.a(n9465), .b(n9464), .O(n9466));
  invx  g08594(.a(n7890), .O(n9467));
  andx  g08595(.a(n7897), .b(n9467), .O(n9468));
  andx  g08596(.a(n7896), .b(n7890), .O(n9469));
  orx   g08597(.a(n9469), .b(n9468), .O(n9470));
  andx  g08598(.a(n9470), .b(n1790), .O(n9471));
  andx  g08599(.a(n9471), .b(n9466), .O(n9472));
  andx  g08600(.a(n7907), .b(n1790), .O(n9473));
  andx  g08601(.a(n9395), .b(n9392), .O(n9474));
  andx  g08602(.a(n9446), .b(n9444), .O(n9475));
  orx   g08603(.a(n9475), .b(n9474), .O(n9476));
  andx  g08604(.a(n9476), .b(n9432), .O(n9477));
  invx  g08605(.a(n9477), .O(n9478));
  orx   g08606(.a(n9476), .b(n9432), .O(n9479));
  andx  g08607(.a(n9479), .b(n9478), .O(n9480));
  andx  g08608(.a(n9480), .b(n9473), .O(n9481));
  andx  g08609(.a(n8351), .b(n1790), .O(n9482));
  andx  g08610(.a(n9377), .b(n9374), .O(n9483));
  andx  g08611(.a(n9438), .b(n9373), .O(n9484));
  orx   g08612(.a(n9484), .b(n9483), .O(n9485));
  andx  g08613(.a(n9485), .b(n9436), .O(n9486));
  invx  g08614(.a(n9486), .O(n9487));
  orx   g08615(.a(n9485), .b(n9436), .O(n9488));
  andx  g08616(.a(n9488), .b(n9487), .O(n9489));
  andx  g08617(.a(n9489), .b(n9482), .O(n9490));
  andx  g08618(.a(n9355), .b(n9350), .O(n9491));
  andx  g08619(.a(n9356), .b(n9349), .O(n9492));
  orx   g08620(.a(n9492), .b(n9491), .O(n9493));
  andx  g08621(.a(n9493), .b(n9353), .O(n9494));
  invx  g08622(.a(n9494), .O(n9495));
  orx   g08623(.a(n9493), .b(n9353), .O(n9496));
  andx  g08624(.a(n9496), .b(n9495), .O(n9497));
  andx  g08625(.a(n8131), .b(n1790), .O(n9498));
  andx  g08626(.a(n9498), .b(n9497), .O(n9499));
  andx  g08627(.a(n9347), .b(n9342), .O(n9500));
  andx  g08628(.a(n9346), .b(n9341), .O(n9501));
  orx   g08629(.a(n9501), .b(n9500), .O(n9502));
  andx  g08630(.a(n9502), .b(n9311), .O(n9503));
  invx  g08631(.a(n9503), .O(n9504));
  orx   g08632(.a(n9502), .b(n9311), .O(n9505));
  andx  g08633(.a(n9505), .b(n9504), .O(n9506));
  andx  g08634(.a(n9338), .b(n9336), .O(n9507));
  andx  g08635(.a(n9339), .b(n9332), .O(n9508));
  orx   g08636(.a(n9508), .b(n9507), .O(n9509));
  andx  g08637(.a(n9509), .b(n9322), .O(n9510));
  invx  g08638(.a(n9510), .O(n9511));
  orx   g08639(.a(n9509), .b(n9322), .O(n9512));
  andx  g08640(.a(n9512), .b(n9511), .O(n9513));
  invx  g08641(.a(n9513), .O(n9514));
  andx  g08642(.a(n7982), .b(n1790), .O(n9515));
  invx  g08643(.a(n9515), .O(n9516));
  andx  g08644(.a(n9516), .b(n9514), .O(n9517));
  invx  g08645(.a(n9517), .O(n9518));
  andx  g08646(.a(n9515), .b(n9513), .O(n9519));
  invx  g08647(.a(n9326), .O(n9520));
  andx  g08648(.a(n9330), .b(n9520), .O(n9521));
  invx  g08649(.a(n9521), .O(n9522));
  andx  g08650(.a(n9522), .b(n9328), .O(n9523));
  invx  g08651(.a(n9523), .O(n9524));
  orx   g08652(.a(n9522), .b(n9328), .O(n9525));
  andx  g08653(.a(n9525), .b(n9524), .O(n9526));
  invx  g08654(.a(n9526), .O(n9527));
  andx  g08655(.a(n7924), .b(n1790), .O(n9528));
  andx  g08656(.a(n9528), .b(n9527), .O(n9529));
  andx  g08657(.a(n9526), .b(n8009), .O(n9530));
  invx  g08658(.a(n9530), .O(n9531));
  invx  g08659(.a(n9323), .O(n9532));
  andx  g08660(.a(n7791), .b(n3230), .O(n9533));
  andx  g08661(.a(n9533), .b(n9532), .O(n9534));
  invx  g08662(.a(n9534), .O(n9535));
  orx   g08663(.a(n9533), .b(n9532), .O(n9536));
  andx  g08664(.a(n9536), .b(n9535), .O(n9537));
  invx  g08665(.a(n9537), .O(n9538));
  andx  g08666(.a(n9538), .b(n9324), .O(n9539));
  andx  g08667(.a(n9324), .b(n7931), .O(n9540));
  andx  g08668(.a(n9538), .b(n7931), .O(n9541));
  orx   g08669(.a(n9541), .b(n9540), .O(n9542));
  orx   g08670(.a(n9542), .b(n9539), .O(n9543));
  andx  g08671(.a(n9543), .b(n1790), .O(n9544));
  andx  g08672(.a(n9544), .b(n9531), .O(n9545));
  orx   g08673(.a(n9545), .b(n9529), .O(n9546));
  orx   g08674(.a(n9546), .b(n9519), .O(n9547));
  andx  g08675(.a(n9547), .b(n9518), .O(n9548));
  andx  g08676(.a(n9548), .b(n9506), .O(n9549));
  orx   g08677(.a(n9548), .b(n9506), .O(n9550));
  andx  g08678(.a(n8062), .b(n1790), .O(n9551));
  andx  g08679(.a(n9551), .b(n9550), .O(n9552));
  orx   g08680(.a(n9552), .b(n9549), .O(n9553));
  andx  g08681(.a(n9553), .b(n9497), .O(n9554));
  andx  g08682(.a(n9553), .b(n9498), .O(n9555));
  orx   g08683(.a(n9555), .b(n9554), .O(n9556));
  orx   g08684(.a(n9556), .b(n9499), .O(n9557));
  orx   g08685(.a(n9371), .b(n9360), .O(n9558));
  andx  g08686(.a(n9558), .b(n9368), .O(n9559));
  invx  g08687(.a(n9559), .O(n9560));
  orx   g08688(.a(n9558), .b(n9368), .O(n9561));
  andx  g08689(.a(n9561), .b(n9560), .O(n9562));
  andx  g08690(.a(n9562), .b(n9557), .O(n9563));
  orx   g08691(.a(n9562), .b(n9557), .O(n9564));
  andx  g08692(.a(n8220), .b(n1790), .O(n9565));
  andx  g08693(.a(n9565), .b(n9564), .O(n9566));
  orx   g08694(.a(n9566), .b(n9563), .O(n9567));
  andx  g08695(.a(n9567), .b(n9482), .O(n9568));
  andx  g08696(.a(n9567), .b(n9489), .O(n9569));
  orx   g08697(.a(n9569), .b(n9568), .O(n9570));
  orx   g08698(.a(n9570), .b(n9490), .O(n9571));
  andx  g08699(.a(n9390), .b(n9433), .O(n9572));
  orx   g08700(.a(n9572), .b(n9388), .O(n9573));
  andx  g08701(.a(n9572), .b(n9388), .O(n9574));
  invx  g08702(.a(n9574), .O(n9575));
  andx  g08703(.a(n9575), .b(n9573), .O(n9576));
  andx  g08704(.a(n9576), .b(n9571), .O(n9577));
  orx   g08705(.a(n9576), .b(n9571), .O(n9578));
  andx  g08706(.a(n8603), .b(n1790), .O(n9579));
  andx  g08707(.a(n9579), .b(n9578), .O(n9580));
  orx   g08708(.a(n9580), .b(n9577), .O(n9581));
  andx  g08709(.a(n9581), .b(n9473), .O(n9582));
  andx  g08710(.a(n9581), .b(n9480), .O(n9583));
  orx   g08711(.a(n9583), .b(n9582), .O(n9584));
  orx   g08712(.a(n9584), .b(n9481), .O(n9585));
  andx  g08713(.a(n9407), .b(n9428), .O(n9586));
  orx   g08714(.a(n9586), .b(n9405), .O(n9587));
  andx  g08715(.a(n9586), .b(n9405), .O(n9588));
  invx  g08716(.a(n9588), .O(n9589));
  andx  g08717(.a(n9589), .b(n9587), .O(n9590));
  andx  g08718(.a(n9590), .b(n9585), .O(n9591));
  orx   g08719(.a(n9590), .b(n9585), .O(n9592));
  andx  g08720(.a(n8852), .b(n1790), .O(n9593));
  andx  g08721(.a(n9593), .b(n9592), .O(n9594));
  orx   g08722(.a(n9594), .b(n9591), .O(n9595));
  andx  g08723(.a(n9050), .b(n1790), .O(n9596));
  andx  g08724(.a(n9596), .b(n9595), .O(n9597));
  andx  g08725(.a(n9412), .b(n9409), .O(n9598));
  andx  g08726(.a(n9454), .b(n9452), .O(n9599));
  orx   g08727(.a(n9599), .b(n9598), .O(n9600));
  andx  g08728(.a(n9600), .b(n9427), .O(n9601));
  invx  g08729(.a(n9601), .O(n9602));
  orx   g08730(.a(n9600), .b(n9427), .O(n9603));
  andx  g08731(.a(n9603), .b(n9602), .O(n9604));
  orx   g08732(.a(n9604), .b(n9597), .O(n9605));
  invx  g08733(.a(n9591), .O(n9606));
  invx  g08734(.a(n9481), .O(n9607));
  invx  g08735(.a(n9473), .O(n9608));
  invx  g08736(.a(n9577), .O(n9609));
  invx  g08737(.a(n9571), .O(n9610));
  invx  g08738(.a(n9573), .O(n9611));
  orx   g08739(.a(n9574), .b(n9611), .O(n9612));
  andx  g08740(.a(n9612), .b(n9610), .O(n9613));
  invx  g08741(.a(n9579), .O(n9614));
  orx   g08742(.a(n9614), .b(n9613), .O(n9615));
  andx  g08743(.a(n9615), .b(n9609), .O(n9616));
  orx   g08744(.a(n9616), .b(n9608), .O(n9617));
  invx  g08745(.a(n9480), .O(n9618));
  orx   g08746(.a(n9616), .b(n9618), .O(n9619));
  andx  g08747(.a(n9619), .b(n9617), .O(n9620));
  andx  g08748(.a(n9620), .b(n9607), .O(n9621));
  invx  g08749(.a(n9587), .O(n9622));
  orx   g08750(.a(n9588), .b(n9622), .O(n9623));
  andx  g08751(.a(n9623), .b(n9621), .O(n9624));
  invx  g08752(.a(n9593), .O(n9625));
  orx   g08753(.a(n9625), .b(n9624), .O(n9626));
  andx  g08754(.a(n9626), .b(n9606), .O(n9627));
  invx  g08755(.a(n9596), .O(n9628));
  andx  g08756(.a(n9628), .b(n9627), .O(n9629));
  invx  g08757(.a(n9629), .O(n9630));
  andx  g08758(.a(n9630), .b(n9605), .O(n9631));
  andx  g08759(.a(n9458), .b(n9414), .O(n9632));
  andx  g08760(.a(n9417), .b(n9456), .O(n9633));
  orx   g08761(.a(n9633), .b(n9632), .O(n9634));
  andx  g08762(.a(n9634), .b(n9424), .O(n9635));
  invx  g08763(.a(n9635), .O(n9636));
  orx   g08764(.a(n9634), .b(n9424), .O(n9637));
  andx  g08765(.a(n9637), .b(n9636), .O(n9638));
  invx  g08766(.a(n9638), .O(n9639));
  andx  g08767(.a(n9639), .b(n9631), .O(n9640));
  andx  g08768(.a(n9267), .b(n1790), .O(n9641));
  andx  g08769(.a(n9641), .b(n9631), .O(n9642));
  invx  g08770(.a(n9641), .O(n9643));
  orx   g08771(.a(n9643), .b(n9638), .O(n9644));
  invx  g08772(.a(n9644), .O(n9645));
  orx   g08773(.a(n9645), .b(n9642), .O(n9646));
  orx   g08774(.a(n9646), .b(n9640), .O(n9647));
  andx  g08775(.a(n9647), .b(n9466), .O(n9648));
  andx  g08776(.a(n9647), .b(n9471), .O(n9649));
  orx   g08777(.a(n9649), .b(n9648), .O(n9650));
  orx   g08778(.a(n9650), .b(n9472), .O(n9651));
  andx  g08779(.a(n9651), .b(n7903), .O(n9652));
  invx  g08780(.a(n7903), .O(n9653));
  invx  g08781(.a(n9472), .O(n9654));
  invx  g08782(.a(n9466), .O(n9655));
  invx  g08783(.a(n9640), .O(n9656));
  orx   g08784(.a(n9628), .b(n9627), .O(n9657));
  invx  g08785(.a(n9604), .O(n9658));
  andx  g08786(.a(n9658), .b(n9657), .O(n9659));
  orx   g08787(.a(n9629), .b(n9659), .O(n9660));
  orx   g08788(.a(n9643), .b(n9660), .O(n9661));
  andx  g08789(.a(n9644), .b(n9661), .O(n9662));
  andx  g08790(.a(n9662), .b(n9656), .O(n9663));
  orx   g08791(.a(n9663), .b(n9655), .O(n9664));
  invx  g08792(.a(n9471), .O(n9665));
  orx   g08793(.a(n9663), .b(n9665), .O(n9666));
  andx  g08794(.a(n9666), .b(n9664), .O(n9667));
  andx  g08795(.a(n9667), .b(n9654), .O(n9668));
  andx  g08796(.a(n9668), .b(n9653), .O(n9669));
  orx   g08797(.a(n9669), .b(n9652), .O(n9670));
  andx  g08798(.a(n8603), .b(n3180), .O(n9671));
  andx  g08799(.a(n8795), .b(n8794), .O(n9672));
  andx  g08800(.a(n8805), .b(n8794), .O(n9673));
  andx  g08801(.a(n8805), .b(n8795), .O(n9674));
  orx   g08802(.a(n9674), .b(n9673), .O(n9675));
  orx   g08803(.a(n9675), .b(n9672), .O(n9676));
  andx  g08804(.a(n9676), .b(n9671), .O(n9677));
  orx   g08805(.a(n8601), .b(n7850), .O(n9678));
  orx   g08806(.a(n7864), .b(n8349), .O(n9679));
  andx  g08807(.a(n9679), .b(n9678), .O(n9680));
  orx   g08808(.a(n9680), .b(n3183), .O(n9681));
  invx  g08809(.a(n9672), .O(n9682));
  orx   g08810(.a(n8800), .b(n8811), .O(n9683));
  orx   g08811(.a(n8800), .b(n8802), .O(n9684));
  andx  g08812(.a(n9684), .b(n9683), .O(n9685));
  andx  g08813(.a(n9685), .b(n9682), .O(n9686));
  andx  g08814(.a(n9686), .b(n9681), .O(n9687));
  orx   g08815(.a(n9687), .b(n9677), .O(n9688));
  orx   g08816(.a(n8742), .b(n8740), .O(n9689));
  orx   g08817(.a(n8736), .b(n8697), .O(n9690));
  andx  g08818(.a(n9690), .b(n9689), .O(n9691));
  andx  g08819(.a(n8749), .b(n8751), .O(n9692));
  andx  g08820(.a(n8755), .b(n8745), .O(n9693));
  orx   g08821(.a(n9693), .b(n9692), .O(n9694));
  andx  g08822(.a(n9694), .b(n9691), .O(n9695));
  orx   g08823(.a(n8758), .b(n9695), .O(n9700));
  andx  g08824(.a(n9700), .b(n8762), .O(n9701));
  andx  g08825(.a(n9700), .b(n8775), .O(n9702));
  andx  g08826(.a(n8775), .b(n8762), .O(n9703));
  orx   g08827(.a(n9703), .b(n9702), .O(n9704));
  orx   g08828(.a(n9704), .b(n9701), .O(n9705));
  orx   g08829(.a(n8675), .b(n3418), .O(n9706));
  orx   g08830(.a(n9706), .b(n9705), .O(n9707));
  invx  g08831(.a(n9701), .O(n9708));
  orx   g08832(.a(n9694), .b(n9691), .O(n9710));
  andx  g08833(.a(n9710), .b(n8759), .O(n9711));
  orx   g08834(.a(n9711), .b(n8766), .O(n9712));
  orx   g08835(.a(n8766), .b(n8771), .O(n9713));
  andx  g08836(.a(n9713), .b(n9712), .O(n9714));
  andx  g08837(.a(n9714), .b(n9708), .O(n9715));
  andx  g08838(.a(n8220), .b(n3171), .O(n9716));
  orx   g08839(.a(n9716), .b(n9715), .O(n9717));
  andx  g08840(.a(n9717), .b(n9707), .O(n9718));
  andx  g08841(.a(n7982), .b(n3721), .O(n9719));
  invx  g08842(.a(n8710), .O(n9720));
  orx   g08843(.a(n8730), .b(n8728), .O(n9721));
  orx   g08844(.a(n8724), .b(n8718), .O(n9722));
  andx  g08845(.a(n9722), .b(n9721), .O(n9723));
  orx   g08846(.a(n9723), .b(n8705), .O(n9724));
  andx  g08847(.a(n9724), .b(n9720), .O(n9725));
  andx  g08848(.a(n9725), .b(n9719), .O(n9726));
  orx   g08849(.a(n7916), .b(n6829), .O(n9727));
  andx  g08850(.a(n7924), .b(n3721), .O(n9728));
  orx   g08851(.a(n9728), .b(n8709), .O(n9729));
  andx  g08852(.a(n8732), .b(n9729), .O(n9730));
  orx   g08853(.a(n9730), .b(n8710), .O(n9731));
  andx  g08854(.a(n9731), .b(n9727), .O(n9732));
  orx   g08855(.a(n9732), .b(n9726), .O(n9733));
  andx  g08856(.a(n8724), .b(n8716), .O(n9734));
  invx  g08857(.a(n9734), .O(n9735));
  andx  g08858(.a(n8716), .b(n8712), .O(n9736));
  invx  g08859(.a(n9736), .O(n9737));
  orx   g08860(.a(n8730), .b(n8715), .O(n9738));
  andx  g08861(.a(n9738), .b(n9737), .O(n9739));
  andx  g08862(.a(n9739), .b(n9735), .O(n9740));
  andx  g08863(.a(n7924), .b(n4063), .O(n9741));
  invx  g08864(.a(n9741), .O(n9742));
  andx  g08865(.a(n9742), .b(n9740), .O(n9743));
  andx  g08866(.a(n8724), .b(n8712), .O(n9744));
  orx   g08867(.a(n9744), .b(n9736), .O(n9745));
  orx   g08868(.a(n9745), .b(n9734), .O(n9746));
  andx  g08869(.a(n9746), .b(n7924), .O(n9747));
  orx   g08870(.a(n9747), .b(n9743), .O(n9748));
  andx  g08871(.a(n7931), .b(n4114), .O(n9749));
  andx  g08872(.a(n9749), .b(n8723), .O(n9750));
  invx  g08873(.a(n9750), .O(n9751));
  orx   g08874(.a(n9749), .b(n8723), .O(n9752));
  andx  g08875(.a(n9752), .b(n9751), .O(n9753));
  andx  g08876(.a(n2724), .b(n7791), .O(n9757));
  andx  g08877(.a(n2723), .b(n4490), .O(n9758));
  andx  g08878(.a(n7792), .b(n4490), .O(n9759));
  orx   g08879(.a(n9759), .b(n9758), .O(n9760));
  andx  g08880(.a(n9760), .b(n7938), .O(n9761));
  orx   g08881(.a(n9761), .b(n9757), .O(n9762));
  andx  g08882(.a(n9762), .b(n9753), .O(n9763));
  invx  g08883(.a(n9752), .O(n9764));
  orx   g08884(.a(n9764), .b(n9750), .O(n9765));
  invx  g08885(.a(n9762), .O(n9766));
  andx  g08886(.a(n9766), .b(n9765), .O(n9767));
  orx   g08887(.a(n9767), .b(n9763), .O(n9768));
  andx  g08888(.a(n9768), .b(n9748), .O(n9769));
  orx   g08889(.a(n9741), .b(n9746), .O(n9770));
  orx   g08890(.a(n9740), .b(n8009), .O(n9771));
  andx  g08891(.a(n9771), .b(n9770), .O(n9772));
  orx   g08892(.a(n9766), .b(n9765), .O(n9773));
  orx   g08893(.a(n9762), .b(n9753), .O(n9774));
  andx  g08894(.a(n9774), .b(n9773), .O(n9775));
  andx  g08895(.a(n9775), .b(n9772), .O(n9776));
  orx   g08896(.a(n9776), .b(n9769), .O(n9777));
  andx  g08897(.a(n9777), .b(n9733), .O(n9778));
  orx   g08898(.a(n9731), .b(n9727), .O(n9779));
  orx   g08899(.a(n9725), .b(n9719), .O(n9780));
  andx  g08900(.a(n9780), .b(n9779), .O(n9781));
  orx   g08901(.a(n9775), .b(n9772), .O(n9782));
  orx   g08902(.a(n9768), .b(n9748), .O(n9783));
  andx  g08903(.a(n9783), .b(n9782), .O(n9784));
  andx  g08904(.a(n9784), .b(n9781), .O(n9785));
  orx   g08905(.a(n9785), .b(n9778), .O(n9786));
  orx   g08906(.a(n8299), .b(n4509), .O(n9787));
  andx  g08907(.a(n8695), .b(n8683), .O(n9788));
  orx   g08908(.a(n8695), .b(n8683), .O(n9789));
  andx  g08909(.a(n9789), .b(n8736), .O(n9790));
  orx   g08910(.a(n9790), .b(n9788), .O(n9791));
  andx  g08911(.a(n9791), .b(n9787), .O(n9792));
  andx  g08912(.a(n8062), .b(n3645), .O(n9793));
  invx  g08913(.a(n9788), .O(n9794));
  andx  g08914(.a(n8689), .b(n8691), .O(n9795));
  orx   g08915(.a(n9795), .b(n8742), .O(n9796));
  andx  g08916(.a(n9796), .b(n9794), .O(n9797));
  andx  g08917(.a(n9797), .b(n9793), .O(n9798));
  orx   g08918(.a(n9798), .b(n9792), .O(n9799));
  andx  g08919(.a(n9799), .b(n9786), .O(n9800));
  orx   g08920(.a(n9784), .b(n9781), .O(n9801));
  orx   g08921(.a(n9777), .b(n9733), .O(n9802));
  andx  g08922(.a(n9802), .b(n9801), .O(n9803));
  orx   g08923(.a(n9797), .b(n9793), .O(n9804));
  orx   g08924(.a(n9791), .b(n9787), .O(n9805));
  andx  g08925(.a(n9805), .b(n9804), .O(n9806));
  andx  g08926(.a(n9806), .b(n9803), .O(n9807));
  orx   g08927(.a(n9807), .b(n9800), .O(n9808));
  orx   g08928(.a(n8770), .b(n4989), .O(n9809));
  andx  g08929(.a(n8749), .b(n9691), .O(n9810));
  orx   g08930(.a(n8749), .b(n9691), .O(n9811));
  andx  g08931(.a(n9811), .b(n8751), .O(n9812));
  orx   g08932(.a(n9812), .b(n9810), .O(n9813));
  andx  g08933(.a(n9813), .b(n9809), .O(n9814));
  andx  g08934(.a(n8131), .b(n3413), .O(n9815));
  orx   g08935(.a(n8755), .b(n8744), .O(n9816));
  andx  g08936(.a(n8755), .b(n8744), .O(n9817));
  orx   g08937(.a(n9817), .b(n8745), .O(n9818));
  andx  g08938(.a(n9818), .b(n9816), .O(n9819));
  andx  g08939(.a(n9819), .b(n9815), .O(n9820));
  orx   g08940(.a(n9820), .b(n9814), .O(n9821));
  andx  g08941(.a(n9821), .b(n9808), .O(n9822));
  orx   g08942(.a(n9806), .b(n9803), .O(n9823));
  orx   g08943(.a(n9799), .b(n9786), .O(n9824));
  andx  g08944(.a(n9824), .b(n9823), .O(n9825));
  orx   g08945(.a(n9819), .b(n9815), .O(n9826));
  orx   g08946(.a(n9813), .b(n9809), .O(n9827));
  andx  g08947(.a(n9827), .b(n9826), .O(n9828));
  andx  g08948(.a(n9828), .b(n9825), .O(n9829));
  orx   g08949(.a(n9829), .b(n9822), .O(n9830));
  orx   g08950(.a(n9830), .b(n9718), .O(n9831));
  andx  g08951(.a(n9716), .b(n9715), .O(n9832));
  andx  g08952(.a(n9706), .b(n9705), .O(n9833));
  orx   g08953(.a(n9833), .b(n9832), .O(n9834));
  orx   g08954(.a(n9828), .b(n9825), .O(n9835));
  orx   g08955(.a(n9821), .b(n9808), .O(n9836));
  andx  g08956(.a(n9836), .b(n9835), .O(n9837));
  orx   g08957(.a(n9837), .b(n9834), .O(n9838));
  andx  g08958(.a(n9838), .b(n9831), .O(n9839));
  andx  g08959(.a(n8218), .b(n8348), .O(n9840));
  orx   g08960(.a(n9840), .b(n7850), .O(n9841));
  orx   g08961(.a(n9841), .b(n3297), .O(n9842));
  andx  g08962(.a(n8792), .b(n8680), .O(n9843));
  orx   g08963(.a(n8792), .b(n8680), .O(n9844));
  andx  g08964(.a(n9844), .b(n8651), .O(n9845));
  orx   g08965(.a(n9845), .b(n9843), .O(n9846));
  andx  g08966(.a(n9846), .b(n9842), .O(n9847));
  andx  g08967(.a(n8351), .b(n3429), .O(n9848));
  orx   g08968(.a(n8785), .b(n8672), .O(n9849));
  andx  g08969(.a(n8785), .b(n8672), .O(n9850));
  orx   g08970(.a(n9850), .b(n8676), .O(n9851));
  andx  g08971(.a(n9851), .b(n9849), .O(n9852));
  andx  g08972(.a(n9852), .b(n9848), .O(n9853));
  orx   g08973(.a(n9853), .b(n9847), .O(n9854));
  andx  g08974(.a(n9854), .b(n9839), .O(n9855));
  andx  g08975(.a(n9837), .b(n9834), .O(n9856));
  andx  g08976(.a(n9830), .b(n9718), .O(n9857));
  orx   g08977(.a(n9857), .b(n9856), .O(n9858));
  orx   g08978(.a(n9852), .b(n9848), .O(n9859));
  orx   g08979(.a(n9846), .b(n9842), .O(n9860));
  andx  g08980(.a(n9860), .b(n9859), .O(n9861));
  andx  g08981(.a(n9861), .b(n9858), .O(n9862));
  orx   g08982(.a(n9862), .b(n9855), .O(n9863));
  orx   g08983(.a(n9863), .b(n9688), .O(n9864));
  orx   g08984(.a(n9686), .b(n9681), .O(n9865));
  orx   g08985(.a(n9676), .b(n9671), .O(n9866));
  andx  g08986(.a(n9866), .b(n9865), .O(n9867));
  orx   g08987(.a(n9861), .b(n9858), .O(n9868));
  orx   g08988(.a(n9854), .b(n9839), .O(n9869));
  andx  g08989(.a(n9869), .b(n9868), .O(n9870));
  orx   g08990(.a(n9870), .b(n9867), .O(n9871));
  andx  g08991(.a(n9871), .b(n9864), .O(n9872));
  andx  g08992(.a(n7907), .b(n3284), .O(n9873));
  invx  g08993(.a(n9873), .O(n9874));
  andx  g08994(.a(n8814), .b(n8811), .O(n9875));
  andx  g08995(.a(n8807), .b(n8794), .O(n9876));
  orx   g08996(.a(n9876), .b(n9875), .O(n9877));
  andx  g08997(.a(n8823), .b(n9877), .O(n9878));
  invx  g08998(.a(n9878), .O(n9879));
  andx  g08999(.a(n8829), .b(n8816), .O(n9880));
  orx   g09000(.a(n9880), .b(n8818), .O(n9881));
  andx  g09001(.a(n9881), .b(n9879), .O(n9882));
  orx   g09002(.a(n9882), .b(n9874), .O(n9883));
  orx   g09003(.a(n8823), .b(n9877), .O(n9884));
  andx  g09004(.a(n9884), .b(n8817), .O(n9885));
  orx   g09005(.a(n9885), .b(n9878), .O(n9886));
  orx   g09006(.a(n9886), .b(n9873), .O(n9887));
  andx  g09007(.a(n9887), .b(n9883), .O(n9888));
  andx  g09008(.a(n9888), .b(n9872), .O(n9889));
  andx  g09009(.a(n9870), .b(n9867), .O(n9890));
  andx  g09010(.a(n9863), .b(n9688), .O(n9891));
  orx   g09011(.a(n9891), .b(n9890), .O(n9892));
  andx  g09012(.a(n9886), .b(n9873), .O(n9893));
  andx  g09013(.a(n9882), .b(n9874), .O(n9894));
  orx   g09014(.a(n9894), .b(n9893), .O(n9895));
  andx  g09015(.a(n9895), .b(n9892), .O(n9896));
  orx   g09016(.a(n9896), .b(n9889), .O(n9897));
  andx  g09017(.a(n8852), .b(n3210), .O(n9898));
  invx  g09018(.a(n9898), .O(n9899));
  orx   g09019(.a(n8831), .b(n9877), .O(n9903));
  andx  g09020(.a(n8823), .b(n8817), .O(n9904));
  andx  g09021(.a(n8829), .b(n8818), .O(n9905));
  orx   g09022(.a(n9905), .b(n9904), .O(n9906));
  orx   g09023(.a(n9906), .b(n8816), .O(n9907));
  andx  g09024(.a(n9907), .b(n9903), .O(n9908));
  andx  g09025(.a(n9908), .b(n7908), .O(n9909));
  andx  g09026(.a(n9908), .b(n8606), .O(n9910));
  andx  g09027(.a(n8606), .b(n7908), .O(n9911));
  orx   g09028(.a(n9911), .b(n9910), .O(n9912));
  orx   g09029(.a(n9912), .b(n9909), .O(n9913));
  andx  g09030(.a(n9913), .b(n9899), .O(n9914));
  invx  g09031(.a(n9909), .O(n9915));
  andx  g09032(.a(n9906), .b(n8816), .O(n9916));
  andx  g09033(.a(n8831), .b(n9877), .O(n9917));
  orx   g09034(.a(n9917), .b(n9916), .O(n9918));
  orx   g09035(.a(n9918), .b(n8648), .O(n9919));
  orx   g09036(.a(n8648), .b(n7909), .O(n9920));
  andx  g09037(.a(n9920), .b(n9919), .O(n9921));
  andx  g09038(.a(n9921), .b(n9915), .O(n9922));
  andx  g09039(.a(n9922), .b(n9898), .O(n9923));
  orx   g09040(.a(n9923), .b(n9914), .O(n9924));
  andx  g09041(.a(n9924), .b(n9897), .O(n9925));
  orx   g09042(.a(n9895), .b(n9892), .O(n9926));
  orx   g09043(.a(n9888), .b(n9872), .O(n9927));
  andx  g09044(.a(n9927), .b(n9926), .O(n9928));
  orx   g09045(.a(n9922), .b(n9898), .O(n9929));
  orx   g09046(.a(n9913), .b(n9899), .O(n9930));
  andx  g09047(.a(n9930), .b(n9929), .O(n9931));
  andx  g09048(.a(n9931), .b(n9928), .O(n9932));
  orx   g09049(.a(n9932), .b(n9925), .O(n9933));
  andx  g09050(.a(n9050), .b(n3221), .O(n9934));
  invx  g09051(.a(n9934), .O(n9935));
  andx  g09052(.a(n9033), .b(n8842), .O(n9936));
  invx  g09053(.a(n9936), .O(n9937));
  andx  g09054(.a(n9024), .b(n9039), .O(n9938));
  orx   g09055(.a(n9938), .b(n9026), .O(n9939));
  andx  g09056(.a(n9939), .b(n9937), .O(n9940));
  orx   g09057(.a(n9940), .b(n9935), .O(n9941));
  orx   g09058(.a(n9033), .b(n8842), .O(n9942));
  andx  g09059(.a(n9942), .b(n8853), .O(n9943));
  orx   g09060(.a(n9943), .b(n9936), .O(n9944));
  orx   g09061(.a(n9944), .b(n9934), .O(n9945));
  andx  g09062(.a(n9945), .b(n9941), .O(n9946));
  andx  g09063(.a(n9946), .b(n9933), .O(n9947));
  orx   g09064(.a(n9931), .b(n9928), .O(n9948));
  orx   g09065(.a(n9924), .b(n9897), .O(n9949));
  andx  g09066(.a(n9949), .b(n9948), .O(n9950));
  andx  g09067(.a(n9944), .b(n9934), .O(n9951));
  andx  g09068(.a(n9940), .b(n9935), .O(n9952));
  orx   g09069(.a(n9952), .b(n9951), .O(n9953));
  andx  g09070(.a(n9953), .b(n9950), .O(n9954));
  orx   g09071(.a(n9954), .b(n9947), .O(n9955));
  andx  g09072(.a(n9267), .b(n3230), .O(n9956));
  invx  g09073(.a(n9956), .O(n9957));
  andx  g09074(.a(n9042), .b(n9039), .O(n9958));
  andx  g09075(.a(n9035), .b(n8842), .O(n9959));
  orx   g09076(.a(n9959), .b(n9958), .O(n9960));
  andx  g09077(.a(n9201), .b(n9960), .O(n9961));
  invx  g09078(.a(n9961), .O(n9962));
  andx  g09079(.a(n9256), .b(n9044), .O(n9963));
  orx   g09080(.a(n9963), .b(n9052), .O(n9964));
  andx  g09081(.a(n9964), .b(n9962), .O(n9965));
  orx   g09082(.a(n9965), .b(n9957), .O(n9966));
  orx   g09083(.a(n9201), .b(n9960), .O(n9967));
  andx  g09084(.a(n9967), .b(n9051), .O(n9968));
  orx   g09085(.a(n9968), .b(n9961), .O(n9969));
  orx   g09086(.a(n9969), .b(n9956), .O(n9970));
  andx  g09087(.a(n9970), .b(n9966), .O(n9971));
  andx  g09088(.a(n9971), .b(n9955), .O(n9972));
  orx   g09089(.a(n9953), .b(n9950), .O(n9973));
  orx   g09090(.a(n9946), .b(n9933), .O(n9974));
  andx  g09091(.a(n9974), .b(n9973), .O(n9975));
  andx  g09092(.a(n9969), .b(n9956), .O(n9976));
  andx  g09093(.a(n9965), .b(n9957), .O(n9977));
  orx   g09094(.a(n9977), .b(n9976), .O(n9978));
  andx  g09095(.a(n9978), .b(n9975), .O(n9979));
  orx   g09096(.a(n9979), .b(n9972), .O(n9980));
  andx  g09097(.a(n9470), .b(n3258), .O(n9981));
  invx  g09098(.a(n9261), .O(n9982));
  orx   g09099(.a(n9982), .b(n9259), .O(n9983));
  andx  g09100(.a(n9419), .b(n9983), .O(n9984));
  orx   g09101(.a(n9419), .b(n9983), .O(n9985));
  andx  g09102(.a(n9985), .b(n9268), .O(n9986));
  orx   g09103(.a(n9986), .b(n9984), .O(n9987));
  andx  g09104(.a(n9987), .b(n9981), .O(n9988));
  invx  g09105(.a(n9981), .O(n9989));
  invx  g09106(.a(n9984), .O(n9990));
  andx  g09107(.a(n9460), .b(n9262), .O(n9991));
  orx   g09108(.a(n9991), .b(n9421), .O(n9992));
  andx  g09109(.a(n9992), .b(n9990), .O(n9993));
  andx  g09110(.a(n9993), .b(n9989), .O(n9994));
  orx   g09111(.a(n9994), .b(n9988), .O(n9995));
  invx  g09112(.a(n9995), .O(n9996));
  andx  g09113(.a(n9996), .b(n9980), .O(n9997));
  orx   g09114(.a(n9978), .b(n9975), .O(n9998));
  orx   g09115(.a(n9971), .b(n9955), .O(n9999));
  andx  g09116(.a(n9999), .b(n9998), .O(n10000));
  andx  g09117(.a(n9995), .b(n10000), .O(n10001));
  orx   g09118(.a(n10001), .b(n9997), .O(n10002));
  orx   g09119(.a(n10002), .b(n9670), .O(n10003));
  invx  g09120(.a(n9670), .O(n10004));
  invx  g09121(.a(n10002), .O(n10005));
  orx   g09122(.a(n10005), .b(n10004), .O(n10006));
  andx  g09123(.a(n10006), .b(n10003), .O(po05));
  andx  g09124(.a(n7982), .b(n4063), .O(n10008));
  orx   g09125(.a(n9775), .b(n9743), .O(n10009));
  andx  g09126(.a(n10009), .b(n9771), .O(n10010));
  orx   g09127(.a(n10010), .b(n10008), .O(n10011));
  orx   g09128(.a(n7916), .b(n4062), .O(n10012));
  andx  g09129(.a(n9768), .b(n9770), .O(n10013));
  orx   g09130(.a(n10013), .b(n9747), .O(n10014));
  orx   g09131(.a(n10014), .b(n10012), .O(n10015));
  andx  g09132(.a(n10015), .b(n10011), .O(n10016));
  andx  g09133(.a(n7938), .b(n2724), .O(n10017));
  andx  g09134(.a(n10017), .b(n8719), .O(n10024));
  andx  g09135(.a(n9762), .b(n9749), .O(n10033));
  orx   g09136(.a(n10033), .b(n8722), .O(n10034));
  andx  g09137(.a(n7924), .b(n4114), .O(n10036));
  orx   g09138(.a(n10036), .b(n10034), .O(n10037));
  andx  g09139(.a(n10034), .b(n7924), .O(n10038));
  invx  g09140(.a(n10038), .O(n10039));
  andx  g09141(.a(n10039), .b(n10037), .O(n10040));
  andx  g09142(.a(n10040), .b(n7959), .O(n10041));
  invx  g09143(.a(n10037), .O(n10042));
  orx   g09144(.a(n10038), .b(n10042), .O(n10043));
  andx  g09145(.a(n10043), .b(n7931), .O(n10044));
  orx   g09146(.a(n10044), .b(n10041), .O(n10045));
  orx   g09147(.a(n10045), .b(n10016), .O(n10046));
  andx  g09148(.a(n10014), .b(n10012), .O(n10047));
  andx  g09149(.a(n10010), .b(n10008), .O(n10048));
  orx   g09150(.a(n10048), .b(n10047), .O(n10049));
  orx   g09151(.a(n10043), .b(n7931), .O(n10050));
  orx   g09152(.a(n10040), .b(n7959), .O(n10051));
  andx  g09153(.a(n10051), .b(n10050), .O(n10052));
  orx   g09154(.a(n10052), .b(n10049), .O(n10053));
  andx  g09155(.a(n10053), .b(n10046), .O(n10054));
  orx   g09156(.a(n8299), .b(n6829), .O(n10055));
  andx  g09157(.a(n9731), .b(n9719), .O(n10056));
  orx   g09158(.a(n9731), .b(n9719), .O(n10057));
  andx  g09159(.a(n10057), .b(n9777), .O(n10058));
  orx   g09160(.a(n10058), .b(n10056), .O(n10059));
  andx  g09161(.a(n10059), .b(n10055), .O(n10060));
  andx  g09162(.a(n8062), .b(n3721), .O(n10061));
  invx  g09163(.a(n10056), .O(n10062));
  andx  g09164(.a(n9725), .b(n9727), .O(n10063));
  orx   g09165(.a(n10063), .b(n9784), .O(n10064));
  andx  g09166(.a(n10064), .b(n10062), .O(n10065));
  andx  g09167(.a(n10065), .b(n10061), .O(n10066));
  orx   g09168(.a(n10066), .b(n10060), .O(n10067));
  andx  g09169(.a(n8131), .b(n3645), .O(n10072));
  orx   g09170(.a(n9797), .b(n9786), .O(n10073));
  andx  g09171(.a(n9797), .b(n9786), .O(n10074));
  orx   g09172(.a(n10074), .b(n9787), .O(n10075));
  andx  g09173(.a(n10075), .b(n10073), .O(n10076));
  orx   g09174(.a(n10076), .b(n10072), .O(n10077));
  orx   g09175(.a(n8770), .b(n4509), .O(n10078));
  andx  g09176(.a(n9791), .b(n9803), .O(n10079));
  orx   g09177(.a(n9791), .b(n9803), .O(n10080));
  andx  g09178(.a(n10080), .b(n9793), .O(n10081));
  orx   g09179(.a(n10081), .b(n10079), .O(n10082));
  orx   g09180(.a(n10082), .b(n10078), .O(n10083));
  andx  g09181(.a(n10083), .b(n10077), .O(n10084));
  orx   g09182(.a(n10084), .b(n10500), .O(n10085));
  andx  g09183(.a(n10082), .b(n10078), .O(n10088));
  andx  g09184(.a(n10076), .b(n10072), .O(n10089));
  orx   g09185(.a(n10089), .b(n10088), .O(n10090));
  orx   g09186(.a(n10090), .b(n10505), .O(n10091));
  andx  g09187(.a(n10091), .b(n10085), .O(n10092));
  andx  g09188(.a(n9815), .b(n9808), .O(n10093));
  orx   g09189(.a(n9815), .b(n9808), .O(n10094));
  andx  g09190(.a(n10094), .b(n9813), .O(n10095));
  orx   g09191(.a(n10095), .b(n10093), .O(n10096));
  orx   g09192(.a(n8675), .b(n4989), .O(n10097));
  orx   g09193(.a(n10097), .b(n10096), .O(n10098));
  invx  g09194(.a(n10093), .O(n10099));
  andx  g09195(.a(n9809), .b(n9825), .O(n10100));
  orx   g09196(.a(n10100), .b(n9819), .O(n10101));
  andx  g09197(.a(n10101), .b(n10099), .O(n10102));
  andx  g09198(.a(n8220), .b(n3413), .O(n10103));
  orx   g09199(.a(n10103), .b(n10102), .O(n10104));
  andx  g09200(.a(n10104), .b(n10098), .O(n10105));
  andx  g09201(.a(n10105), .b(n10092), .O(n10106));
  andx  g09202(.a(n10090), .b(n10505), .O(n10107));
  andx  g09203(.a(n10084), .b(n10500), .O(n10108));
  orx   g09204(.a(n10108), .b(n10107), .O(n10109));
  andx  g09205(.a(n10103), .b(n10102), .O(n10110));
  andx  g09206(.a(n10097), .b(n10096), .O(n10111));
  orx   g09207(.a(n10111), .b(n10110), .O(n10112));
  andx  g09208(.a(n10112), .b(n10109), .O(n10113));
  orx   g09209(.a(n10113), .b(n10106), .O(n10114));
  orx   g09210(.a(n9841), .b(n3418), .O(n10115));
  andx  g09211(.a(n9837), .b(n9705), .O(n10116));
  orx   g09212(.a(n9837), .b(n9705), .O(n10117));
  andx  g09213(.a(n10117), .b(n9716), .O(n10118));
  orx   g09214(.a(n10118), .b(n10116), .O(n10119));
  andx  g09215(.a(n10119), .b(n10115), .O(n10120));
  andx  g09216(.a(n8351), .b(n3171), .O(n10121));
  orx   g09217(.a(n9830), .b(n9715), .O(n10122));
  andx  g09218(.a(n9830), .b(n9715), .O(n10123));
  orx   g09219(.a(n10123), .b(n9706), .O(n10124));
  andx  g09220(.a(n10124), .b(n10122), .O(n10125));
  andx  g09221(.a(n10125), .b(n10121), .O(n10126));
  orx   g09222(.a(n10126), .b(n10120), .O(n10127));
  andx  g09223(.a(n10127), .b(n10114), .O(n10128));
  orx   g09224(.a(n10112), .b(n10109), .O(n10129));
  orx   g09225(.a(n10105), .b(n10092), .O(n10130));
  andx  g09226(.a(n10130), .b(n10129), .O(n10131));
  orx   g09227(.a(n10125), .b(n10121), .O(n10132));
  orx   g09228(.a(n10119), .b(n10115), .O(n10133));
  andx  g09229(.a(n10133), .b(n10132), .O(n10134));
  andx  g09230(.a(n10134), .b(n10131), .O(n10135));
  orx   g09231(.a(n10135), .b(n10128), .O(n10136));
  andx  g09232(.a(n8603), .b(n3429), .O(n10137));
  andx  g09233(.a(n9848), .b(n9839), .O(n10138));
  orx   g09234(.a(n9848), .b(n9839), .O(n10139));
  andx  g09235(.a(n10139), .b(n9846), .O(n10140));
  orx   g09236(.a(n10140), .b(n10138), .O(n10141));
  andx  g09237(.a(n10141), .b(n10137), .O(n10142));
  orx   g09238(.a(n9680), .b(n3297), .O(n10143));
  invx  g09239(.a(n10138), .O(n10144));
  andx  g09240(.a(n9842), .b(n9858), .O(n10145));
  orx   g09241(.a(n10145), .b(n9852), .O(n10146));
  andx  g09242(.a(n10146), .b(n10144), .O(n10147));
  andx  g09243(.a(n10147), .b(n10143), .O(n10148));
  orx   g09244(.a(n10148), .b(n10142), .O(n10149));
  orx   g09245(.a(n10149), .b(n10136), .O(n10150));
  andx  g09246(.a(n10149), .b(n10136), .O(n10152));
  andx  g09247(.a(n7907), .b(n3180), .O(n10154));
  orx   g09248(.a(n9863), .b(n9686), .O(n10155));
  andx  g09249(.a(n9863), .b(n9686), .O(n10156));
  orx   g09250(.a(n10156), .b(n9681), .O(n10157));
  andx  g09251(.a(n10157), .b(n10155), .O(n10158));
  orx   g09252(.a(n10158), .b(n10154), .O(n10159));
  invx  g09253(.a(n7906), .O(n10160));
  andx  g09254(.a(n10160), .b(n7904), .O(n10161));
  orx   g09255(.a(n10161), .b(n3183), .O(n10162));
  andx  g09256(.a(n9870), .b(n9676), .O(n10163));
  orx   g09257(.a(n9870), .b(n9676), .O(n10164));
  andx  g09258(.a(n10164), .b(n9671), .O(n10165));
  orx   g09259(.a(n10165), .b(n10163), .O(n10166));
  orx   g09260(.a(n10166), .b(n10162), .O(n10167));
  andx  g09261(.a(n10167), .b(n10159), .O(n10168));
  orx   g09262(.a(n10168), .b(n10383), .O(n10169));
  andx  g09263(.a(n10166), .b(n10162), .O(n10172));
  andx  g09264(.a(n10158), .b(n10154), .O(n10173));
  orx   g09265(.a(n10173), .b(n10172), .O(n10174));
  orx   g09266(.a(n10174), .b(n10388), .O(n10175));
  andx  g09267(.a(n10175), .b(n10169), .O(n10176));
  andx  g09268(.a(n8852), .b(n3284), .O(n10177));
  invx  g09269(.a(n10177), .O(n10178));
  andx  g09270(.a(n9873), .b(n9872), .O(n10179));
  orx   g09271(.a(n9873), .b(n9872), .O(n10180));
  andx  g09272(.a(n10180), .b(n9886), .O(n10181));
  orx   g09273(.a(n10181), .b(n10179), .O(n10182));
  andx  g09274(.a(n10182), .b(n10178), .O(n10183));
  invx  g09275(.a(n10179), .O(n10184));
  andx  g09276(.a(n9874), .b(n9892), .O(n10185));
  orx   g09277(.a(n10185), .b(n9882), .O(n10186));
  andx  g09278(.a(n10186), .b(n10184), .O(n10187));
  andx  g09279(.a(n10187), .b(n10177), .O(n10188));
  orx   g09280(.a(n10188), .b(n10183), .O(n10189));
  andx  g09281(.a(n10189), .b(n10176), .O(n10190));
  andx  g09282(.a(n10174), .b(n10388), .O(n10191));
  andx  g09283(.a(n10168), .b(n10383), .O(n10192));
  orx   g09284(.a(n10192), .b(n10191), .O(n10193));
  orx   g09285(.a(n10187), .b(n10177), .O(n10194));
  orx   g09286(.a(n10182), .b(n10178), .O(n10195));
  andx  g09287(.a(n10195), .b(n10194), .O(n10196));
  andx  g09288(.a(n10196), .b(n10193), .O(n10197));
  orx   g09289(.a(n10197), .b(n10190), .O(n10198));
  andx  g09290(.a(n9050), .b(n3210), .O(n10199));
  andx  g09291(.a(n9913), .b(n9928), .O(n10200));
  invx  g09292(.a(n10200), .O(n10201));
  andx  g09293(.a(n9922), .b(n9897), .O(n10202));
  orx   g09294(.a(n10202), .b(n9899), .O(n10203));
  andx  g09295(.a(n10203), .b(n10201), .O(n10204));
  orx   g09296(.a(n10204), .b(n10199), .O(n10205));
  invx  g09297(.a(n10199), .O(n10206));
  orx   g09298(.a(n9913), .b(n9928), .O(n10207));
  andx  g09299(.a(n10207), .b(n9898), .O(n10208));
  orx   g09300(.a(n10208), .b(n10200), .O(n10209));
  orx   g09301(.a(n10209), .b(n10206), .O(n10210));
  andx  g09302(.a(n10210), .b(n10205), .O(n10211));
  orx   g09303(.a(n10211), .b(n10198), .O(n10212));
  orx   g09304(.a(n10196), .b(n10193), .O(n10213));
  orx   g09305(.a(n10189), .b(n10176), .O(n10214));
  andx  g09306(.a(n10214), .b(n10213), .O(n10215));
  andx  g09307(.a(n10209), .b(n10206), .O(n10216));
  andx  g09308(.a(n10204), .b(n10199), .O(n10217));
  orx   g09309(.a(n10217), .b(n10216), .O(n10218));
  orx   g09310(.a(n10218), .b(n10215), .O(n10219));
  andx  g09311(.a(n10219), .b(n10212), .O(n10220));
  andx  g09312(.a(n9267), .b(n3221), .O(n10221));
  invx  g09313(.a(n10221), .O(n10222));
  andx  g09314(.a(n9934), .b(n9933), .O(n10223));
  orx   g09315(.a(n9934), .b(n9933), .O(n10224));
  andx  g09316(.a(n10224), .b(n9944), .O(n10225));
  orx   g09317(.a(n10225), .b(n10223), .O(n10226));
  andx  g09318(.a(n10226), .b(n10222), .O(n10227));
  invx  g09319(.a(n10223), .O(n10228));
  andx  g09320(.a(n9935), .b(n9950), .O(n10229));
  orx   g09321(.a(n10229), .b(n9940), .O(n10230));
  andx  g09322(.a(n10230), .b(n10228), .O(n10231));
  andx  g09323(.a(n10231), .b(n10221), .O(n10232));
  orx   g09324(.a(n10232), .b(n10227), .O(n10233));
  andx  g09325(.a(n10233), .b(n10220), .O(n10234));
  andx  g09326(.a(n10218), .b(n10215), .O(n10235));
  andx  g09327(.a(n10211), .b(n10198), .O(n10236));
  orx   g09328(.a(n10236), .b(n10235), .O(n10237));
  orx   g09329(.a(n10231), .b(n10221), .O(n10238));
  orx   g09330(.a(n10226), .b(n10222), .O(n10239));
  andx  g09331(.a(n10239), .b(n10238), .O(n10240));
  andx  g09332(.a(n10240), .b(n10237), .O(n10241));
  orx   g09333(.a(n10241), .b(n10234), .O(n10242));
  andx  g09334(.a(n9969), .b(n9975), .O(n10243));
  invx  g09335(.a(n10243), .O(n10244));
  andx  g09336(.a(n9965), .b(n9955), .O(n10245));
  orx   g09337(.a(n10245), .b(n9957), .O(n10246));
  andx  g09338(.a(n10246), .b(n10244), .O(n10247));
  andx  g09339(.a(n9470), .b(n3230), .O(n10248));
  invx  g09340(.a(n10248), .O(n10249));
  andx  g09341(.a(n10249), .b(n10247), .O(n10250));
  orx   g09342(.a(n9969), .b(n9975), .O(n10251));
  andx  g09343(.a(n10251), .b(n9956), .O(n10252));
  orx   g09344(.a(n10252), .b(n10243), .O(n10253));
  andx  g09345(.a(n10248), .b(n10253), .O(n10254));
  orx   g09346(.a(n10254), .b(n10250), .O(n10255));
  orx   g09347(.a(n10255), .b(n10242), .O(n10256));
  orx   g09348(.a(n10240), .b(n10237), .O(n10257));
  orx   g09349(.a(n10233), .b(n10220), .O(n10258));
  andx  g09350(.a(n10258), .b(n10257), .O(n10259));
  orx   g09351(.a(n10248), .b(n10253), .O(n10260));
  orx   g09352(.a(n10249), .b(n10247), .O(n10261));
  andx  g09353(.a(n10261), .b(n10260), .O(n10262));
  orx   g09354(.a(n10262), .b(n10259), .O(n10263));
  andx  g09355(.a(n10263), .b(n10256), .O(n10264));
  andx  g09356(.a(n7902), .b(n3258), .O(n10265));
  invx  g09357(.a(n10265), .O(n10266));
  andx  g09358(.a(n9981), .b(n9980), .O(n10267));
  orx   g09359(.a(n9981), .b(n9980), .O(n10268));
  andx  g09360(.a(n10268), .b(n9987), .O(n10269));
  orx   g09361(.a(n10269), .b(n10267), .O(n10270));
  andx  g09362(.a(n10270), .b(n10266), .O(n10271));
  invx  g09363(.a(n10267), .O(n10272));
  andx  g09364(.a(n9989), .b(n10000), .O(n10273));
  orx   g09365(.a(n10273), .b(n9993), .O(n10274));
  andx  g09366(.a(n10274), .b(n10272), .O(n10275));
  andx  g09367(.a(n10275), .b(n10265), .O(n10276));
  orx   g09368(.a(n10276), .b(n10271), .O(n10277));
  andx  g09369(.a(n10277), .b(n10264), .O(n10278));
  invx  g09370(.a(n10278), .O(n10279));
  orx   g09371(.a(n10277), .b(n10264), .O(n10280));
  andx  g09372(.a(n10280), .b(n10279), .O(n10281));
  andx  g09373(.a(n10005), .b(n9651), .O(n10282));
  invx  g09374(.a(n10282), .O(n10283));
  andx  g09375(.a(n10002), .b(n9668), .O(n10284));
  orx   g09376(.a(n10284), .b(n9653), .O(n10285));
  andx  g09377(.a(n10285), .b(n10283), .O(n10286));
  andx  g09378(.a(n7898), .b(n7732), .O(n10287));
  invx  g09379(.a(n10287), .O(n10288));
  andx  g09380(.a(n7659), .b(n7657), .O(n10289));
  orx   g09381(.a(n10289), .b(n7727), .O(n10290));
  andx  g09382(.a(n7689), .b(n7669), .O(n10293));
  invx  g09383(.a(n10293), .O(n10294));
  andx  g09384(.a(n7691), .b(n7668), .O(n10295));
  orx   g09385(.a(n10295), .b(n7671), .O(n10296));
  andx  g09386(.a(n10296), .b(n10294), .O(n10297));
  invx  g09387(.a(n10297), .O(n10298));
  andx  g09388(.a(n10297), .b(n299), .O(n10300));
  andx  g09389(.a(n4114), .b(n827), .O(n10302));
  invx  g09390(.a(n10302), .O(n10303));
  andx  g09391(.a(n7684), .b(n5799), .O(n10307));
  orx   g09392(.a(n10307), .b(n4062), .O(n10308));
  andx  g09393(.a(n7685), .b(n3721), .O(n10309));
  invx  g09394(.a(n10309), .O(n10310));
  andx  g09395(.a(n10310), .b(n10308), .O(n10311));
  invx  g09396(.a(n10311), .O(n10312));
  andx  g09397(.a(n10312), .b(n4063), .O(n10313));
  invx  g09398(.a(n10313), .O(n10314));
  orx   g09399(.a(n10312), .b(n4063), .O(n10315));
  andx  g09400(.a(n10315), .b(n10314), .O(n10316));
  andx  g09401(.a(n10316), .b(n10300), .O(n10317));
  invx  g09402(.a(n10317), .O(n10318));
  orx   g09403(.a(n10316), .b(n10300), .O(n10319));
  andx  g09404(.a(n10319), .b(n10318), .O(n10320));
  invx  g09405(.a(n10320), .O(n10321));
  andx  g09406(.a(n338), .b(n7703), .O(n10322));
  orx   g09407(.a(n10322), .b(n7695), .O(n10323));
  andx  g09408(.a(n10323), .b(n2724), .O(n10324));
  invx  g09409(.a(n10323), .O(n10329));
  andx  g09410(.a(n10329), .b(n10321), .O(n10330));
  orx   g09411(.a(n10695), .b(n10330), .O(n10332));
  andx  g09412(.a(n7707), .b(n7706), .O(n10333));
  invx  g09413(.a(n10333), .O(n10334));
  orx   g09414(.a(n7705), .b(n7709), .O(n10336));
  andx  g09415(.a(n10336), .b(n10334), .O(n10337));
  andx  g09416(.a(n10337), .b(n10332), .O(n10338));
  orx   g09417(.a(n10337), .b(n10332), .O(n10339));
  invx  g09418(.a(n10339), .O(n10340));
  orx   g09419(.a(n10340), .b(n10338), .O(n10341));
  andx  g09420(.a(n7721), .b(n7661), .O(n10342));
  invx  g09421(.a(n10342), .O(n10343));
  andx  g09422(.a(n10343), .b(n10341), .O(n10344));
  invx  g09423(.a(n10344), .O(n10345));
  orx   g09424(.a(n10343), .b(n10341), .O(n10346));
  andx  g09425(.a(n10346), .b(n10345), .O(n10347));
  invx  g09426(.a(n10347), .O(n10348));
  andx  g09427(.a(n10348), .b(n10290), .O(n10349));
  invx  g09428(.a(n10290), .O(n10350));
  andx  g09429(.a(n10347), .b(n10350), .O(n10351));
  orx   g09430(.a(n10351), .b(n10349), .O(n10352));
  andx  g09431(.a(n10352), .b(n10288), .O(n10353));
  invx  g09432(.a(n10352), .O(n10354));
  andx  g09433(.a(n10354), .b(n10287), .O(n10355));
  orx   g09434(.a(n10355), .b(n10353), .O(n10356));
  andx  g09435(.a(n10356), .b(n1790), .O(n10357));
  invx  g09436(.a(n10357), .O(n10358));
  andx  g09437(.a(n10358), .b(n10286), .O(n10359));
  orx   g09438(.a(n10005), .b(n9651), .O(n10360));
  andx  g09439(.a(n10360), .b(n7903), .O(n10361));
  orx   g09440(.a(n10361), .b(n10282), .O(n10362));
  andx  g09441(.a(n10357), .b(n10362), .O(n10363));
  orx   g09442(.a(n10363), .b(n10359), .O(n10364));
  invx  g09443(.a(n10364), .O(n10365));
  andx  g09444(.a(n10365), .b(n10281), .O(n10366));
  invx  g09445(.a(n10281), .O(n10367));
  andx  g09446(.a(n10364), .b(n10367), .O(n10368));
  orx   g09447(.a(n10368), .b(n10366), .O(po06));
  andx  g09448(.a(n8852), .b(n3180), .O(n10370));
  invx  g09449(.a(n10370), .O(n10371));
  orx   g09450(.a(n10134), .b(n10131), .O(n10376));
  orx   g09451(.a(n10127), .b(n10114), .O(n10377));
  andx  g09452(.a(n10377), .b(n10376), .O(n10378));
  andx  g09453(.a(n10147), .b(n10137), .O(n10379));
  andx  g09454(.a(n10141), .b(n10143), .O(n10380));
  orx   g09455(.a(n10380), .b(n10379), .O(n10381));
  andx  g09456(.a(n10381), .b(n10378), .O(n10382));
  orx   g09457(.a(n10382), .b(n10152), .O(n10383));
  andx  g09458(.a(n10383), .b(n10154), .O(n10384));
  invx  g09459(.a(n10384), .O(n10385));
  orx   g09460(.a(n10381), .b(n10378), .O(n10386));
  andx  g09461(.a(n10150), .b(n10386), .O(n10388));
  orx   g09462(.a(n10388), .b(n10158), .O(n10389));
  orx   g09463(.a(n10158), .b(n10162), .O(n10390));
  andx  g09464(.a(n10390), .b(n10389), .O(n10391));
  andx  g09465(.a(n10391), .b(n10385), .O(n10392));
  orx   g09466(.a(n10392), .b(n10371), .O(n10393));
  andx  g09467(.a(n10383), .b(n10166), .O(n10394));
  andx  g09468(.a(n10166), .b(n10154), .O(n10395));
  orx   g09469(.a(n10395), .b(n10394), .O(n10396));
  orx   g09470(.a(n10396), .b(n10384), .O(n10397));
  orx   g09471(.a(n10397), .b(n10370), .O(n10398));
  andx  g09472(.a(n10398), .b(n10393), .O(n10399));
  andx  g09473(.a(n8603), .b(n3171), .O(n10400));
  andx  g09474(.a(n10121), .b(n10131), .O(n10401));
  andx  g09475(.a(n10119), .b(n10131), .O(n10402));
  andx  g09476(.a(n10119), .b(n10121), .O(n10403));
  orx   g09477(.a(n10403), .b(n10402), .O(n10404));
  orx   g09478(.a(n10404), .b(n10401), .O(n10405));
  andx  g09479(.a(n10405), .b(n10400), .O(n10406));
  orx   g09480(.a(n9680), .b(n3418), .O(n10407));
  invx  g09481(.a(n10401), .O(n10408));
  orx   g09482(.a(n10125), .b(n10114), .O(n10409));
  orx   g09483(.a(n10125), .b(n10115), .O(n10410));
  andx  g09484(.a(n10410), .b(n10409), .O(n10411));
  andx  g09485(.a(n10411), .b(n10408), .O(n10412));
  andx  g09486(.a(n10412), .b(n10407), .O(n10413));
  orx   g09487(.a(n10413), .b(n10406), .O(n10414));
  andx  g09488(.a(n8062), .b(n4063), .O(n10415));
  invx  g09489(.a(n10415), .O(n10416));
  andx  g09490(.a(n10045), .b(n10014), .O(n10417));
  andx  g09491(.a(n10045), .b(n10008), .O(n10418));
  andx  g09492(.a(n10014), .b(n10008), .O(n10419));
  orx   g09493(.a(n10419), .b(n10418), .O(n10420));
  orx   g09494(.a(n10420), .b(n10417), .O(n10421));
  andx  g09495(.a(n10421), .b(n10416), .O(n10422));
  invx  g09496(.a(n10417), .O(n10423));
  orx   g09497(.a(n10052), .b(n10012), .O(n10424));
  invx  g09498(.a(n10419), .O(n10425));
  andx  g09499(.a(n10425), .b(n10424), .O(n10426));
  andx  g09500(.a(n10426), .b(n10423), .O(n10427));
  andx  g09501(.a(n10427), .b(n10415), .O(n10428));
  orx   g09502(.a(n10428), .b(n10422), .O(n10429));
  andx  g09503(.a(n7982), .b(n4114), .O(n10430));
  invx  g09504(.a(n10430), .O(n10431));
  andx  g09505(.a(n10037), .b(n7931), .O(n10432));
  orx   g09506(.a(n10432), .b(n10038), .O(n10433));
  orx   g09507(.a(n10433), .b(n10431), .O(n10434));
  invx  g09508(.a(n10434), .O(n10435));
  andx  g09509(.a(n10433), .b(n10431), .O(n10436));
  orx   g09510(.a(n10436), .b(n10435), .O(n10437));
  andx  g09511(.a(n7931), .b(n10017), .O(n10438));
  orx   g09512(.a(n10438), .b(n10024), .O(n10439));
  invx  g09513(.a(n10439), .O(n10440));
  andx  g09514(.a(n7924), .b(n10437), .O(n10453));
  invx  g09515(.a(n10436), .O(n10454));
  andx  g09516(.a(n10454), .b(n10434), .O(n10455));
  andx  g09517(.a(n8009), .b(n10455), .O(n10456));
  orx   g09518(.a(n10456), .b(n10453), .O(n10457));
  orx   g09519(.a(n10457), .b(n10429), .O(n10458));
  orx   g09520(.a(n10427), .b(n10415), .O(n10459));
  orx   g09521(.a(n10421), .b(n10416), .O(n10460));
  andx  g09522(.a(n10460), .b(n10459), .O(n10461));
  orx   g09523(.a(n8009), .b(n10455), .O(n10462));
  orx   g09524(.a(n7924), .b(n10437), .O(n10463));
  andx  g09525(.a(n10463), .b(n10462), .O(n10464));
  orx   g09526(.a(n10464), .b(n10461), .O(n10465));
  andx  g09527(.a(n10465), .b(n10458), .O(n10466));
  andx  g09528(.a(n10052), .b(n10049), .O(n10467));
  andx  g09529(.a(n10045), .b(n10016), .O(n10468));
  orx   g09530(.a(n10468), .b(n10467), .O(n10469));
  andx  g09531(.a(n10059), .b(n10469), .O(n10470));
  orx   g09532(.a(n10059), .b(n10469), .O(n10471));
  andx  g09533(.a(n10471), .b(n10061), .O(n10472));
  orx   g09534(.a(n10472), .b(n10470), .O(n10473));
  andx  g09535(.a(n8131), .b(n3721), .O(n10474));
  orx   g09536(.a(n10474), .b(n10473), .O(n10475));
  invx  g09537(.a(n10470), .O(n10476));
  andx  g09538(.a(n10065), .b(n10054), .O(n10477));
  orx   g09539(.a(n10477), .b(n10055), .O(n10478));
  andx  g09540(.a(n10478), .b(n10476), .O(n10479));
  invx  g09541(.a(n10474), .O(n10480));
  orx   g09542(.a(n10480), .b(n10479), .O(n10481));
  andx  g09543(.a(n10481), .b(n10475), .O(n10482));
  andx  g09544(.a(n10482), .b(n10466), .O(n10483));
  andx  g09545(.a(n10464), .b(n10461), .O(n10484));
  andx  g09546(.a(n10457), .b(n10429), .O(n10485));
  orx   g09547(.a(n10485), .b(n10484), .O(n10486));
  andx  g09548(.a(n10480), .b(n10479), .O(n10487));
  andx  g09549(.a(n10474), .b(n10473), .O(n10488));
  orx   g09550(.a(n10488), .b(n10487), .O(n10489));
  andx  g09551(.a(n10489), .b(n10486), .O(n10490));
  orx   g09552(.a(n10490), .b(n10483), .O(n10491));
  orx   g09553(.a(n10067), .b(n10469), .O(n10495));
  andx  g09554(.a(n10059), .b(n10061), .O(n10496));
  andx  g09555(.a(n10065), .b(n10055), .O(n10497));
  orx   g09556(.a(n10497), .b(n10496), .O(n10498));
  orx   g09557(.a(n10498), .b(n10054), .O(n10499));
  andx  g09558(.a(n10499), .b(n10495), .O(n10500));
  andx  g09559(.a(n10500), .b(n10072), .O(n10501));
  invx  g09560(.a(n10501), .O(n10502));
  andx  g09561(.a(n10498), .b(n10054), .O(n10503));
  andx  g09562(.a(n10067), .b(n10469), .O(n10504));
  orx   g09563(.a(n10504), .b(n10503), .O(n10505));
  orx   g09564(.a(n10505), .b(n10076), .O(n10506));
  orx   g09565(.a(n10076), .b(n10078), .O(n10507));
  andx  g09566(.a(n10507), .b(n10506), .O(n10508));
  andx  g09567(.a(n10508), .b(n10502), .O(n10509));
  andx  g09568(.a(n8220), .b(n3645), .O(n10510));
  andx  g09569(.a(n10510), .b(n10509), .O(n10511));
  andx  g09570(.a(n10500), .b(n10082), .O(n10512));
  andx  g09571(.a(n10082), .b(n10072), .O(n10513));
  orx   g09572(.a(n10513), .b(n10512), .O(n10514));
  orx   g09573(.a(n10514), .b(n10501), .O(n10515));
  orx   g09574(.a(n8675), .b(n4509), .O(n10516));
  andx  g09575(.a(n10516), .b(n10515), .O(n10517));
  orx   g09576(.a(n10517), .b(n10511), .O(n10518));
  orx   g09577(.a(n10518), .b(n10491), .O(n10519));
  orx   g09578(.a(n10489), .b(n10486), .O(n10520));
  orx   g09579(.a(n10482), .b(n10466), .O(n10521));
  andx  g09580(.a(n10521), .b(n10520), .O(n10522));
  orx   g09581(.a(n10516), .b(n10515), .O(n10523));
  orx   g09582(.a(n10510), .b(n10509), .O(n10524));
  andx  g09583(.a(n10524), .b(n10523), .O(n10525));
  orx   g09584(.a(n10525), .b(n10522), .O(n10526));
  andx  g09585(.a(n10526), .b(n10519), .O(n10527));
  andx  g09586(.a(n8351), .b(n3413), .O(n10528));
  orx   g09587(.a(n10102), .b(n10092), .O(n10529));
  andx  g09588(.a(n10102), .b(n10092), .O(n10530));
  orx   g09589(.a(n10530), .b(n10097), .O(n10531));
  andx  g09590(.a(n10531), .b(n10529), .O(n10532));
  orx   g09591(.a(n10532), .b(n10528), .O(n10533));
  orx   g09592(.a(n9841), .b(n4989), .O(n10534));
  andx  g09593(.a(n10096), .b(n10109), .O(n10535));
  orx   g09594(.a(n10096), .b(n10109), .O(n10536));
  andx  g09595(.a(n10536), .b(n10103), .O(n10537));
  orx   g09596(.a(n10537), .b(n10535), .O(n10538));
  orx   g09597(.a(n10538), .b(n10534), .O(n10539));
  andx  g09598(.a(n10539), .b(n10533), .O(n10540));
  orx   g09599(.a(n10540), .b(n10527), .O(n10541));
  andx  g09600(.a(n10525), .b(n10522), .O(n10542));
  andx  g09601(.a(n10518), .b(n10491), .O(n10543));
  orx   g09602(.a(n10543), .b(n10542), .O(n10544));
  andx  g09603(.a(n10538), .b(n10534), .O(n10545));
  andx  g09604(.a(n10532), .b(n10528), .O(n10546));
  orx   g09605(.a(n10546), .b(n10545), .O(n10547));
  orx   g09606(.a(n10547), .b(n10544), .O(n10548));
  andx  g09607(.a(n10548), .b(n10541), .O(n10549));
  orx   g09608(.a(n10161), .b(n3297), .O(n10554));
  andx  g09609(.a(n10141), .b(n10136), .O(n10555));
  orx   g09610(.a(n10141), .b(n10136), .O(n10556));
  andx  g09611(.a(n10556), .b(n10137), .O(n10557));
  orx   g09612(.a(n10557), .b(n10555), .O(n10558));
  andx  g09613(.a(n10558), .b(n10554), .O(n10559));
  andx  g09614(.a(n7907), .b(n3429), .O(n10560));
  orx   g09615(.a(n10147), .b(n10378), .O(n10561));
  andx  g09616(.a(n10147), .b(n10378), .O(n10562));
  orx   g09617(.a(n10562), .b(n10143), .O(n10563));
  andx  g09618(.a(n10563), .b(n10561), .O(n10564));
  andx  g09619(.a(n10564), .b(n10560), .O(n10565));
  orx   g09620(.a(n10565), .b(n10559), .O(n10566));
  andx  g09621(.a(n10566), .b(n10800), .O(n10567));
  orx   g09622(.a(n10564), .b(n10560), .O(n10570));
  orx   g09623(.a(n10558), .b(n10554), .O(n10571));
  andx  g09624(.a(n10571), .b(n10570), .O(n10572));
  andx  g09625(.a(n10572), .b(n10795), .O(n10573));
  orx   g09626(.a(n10573), .b(n10567), .O(n10574));
  andx  g09627(.a(n10574), .b(n10399), .O(n10575));
  andx  g09628(.a(n10397), .b(n10370), .O(n10576));
  andx  g09629(.a(n10392), .b(n10371), .O(n10577));
  orx   g09630(.a(n10577), .b(n10576), .O(n10578));
  orx   g09631(.a(n10572), .b(n10795), .O(n10579));
  orx   g09632(.a(n10566), .b(n10800), .O(n10580));
  andx  g09633(.a(n10580), .b(n10579), .O(n10581));
  andx  g09634(.a(n10581), .b(n10578), .O(n10582));
  orx   g09635(.a(n10582), .b(n10575), .O(n10583));
  andx  g09636(.a(n8850), .b(n9047), .O(n10584));
  orx   g09637(.a(n10584), .b(n7881), .O(n10585));
  orx   g09638(.a(n10585), .b(n3201), .O(n10586));
  andx  g09639(.a(n10182), .b(n10193), .O(n10587));
  orx   g09640(.a(n10182), .b(n10193), .O(n10588));
  andx  g09641(.a(n10588), .b(n10177), .O(n10589));
  orx   g09642(.a(n10589), .b(n10587), .O(n10590));
  andx  g09643(.a(n10590), .b(n10586), .O(n10591));
  andx  g09644(.a(n9050), .b(n3284), .O(n10592));
  orx   g09645(.a(n10187), .b(n10176), .O(n10593));
  andx  g09646(.a(n10187), .b(n10176), .O(n10594));
  orx   g09647(.a(n10594), .b(n10178), .O(n10595));
  andx  g09648(.a(n10595), .b(n10593), .O(n10596));
  andx  g09649(.a(n10596), .b(n10592), .O(n10597));
  orx   g09650(.a(n10597), .b(n10591), .O(n10598));
  andx  g09651(.a(n10598), .b(n10583), .O(n10599));
  orx   g09652(.a(n10581), .b(n10578), .O(n10600));
  orx   g09653(.a(n10574), .b(n10399), .O(n10601));
  andx  g09654(.a(n10601), .b(n10600), .O(n10602));
  orx   g09655(.a(n10596), .b(n10592), .O(n10603));
  orx   g09656(.a(n10590), .b(n10586), .O(n10604));
  andx  g09657(.a(n10604), .b(n10603), .O(n10605));
  andx  g09658(.a(n10605), .b(n10602), .O(n10606));
  orx   g09659(.a(n10606), .b(n10599), .O(n10607));
  andx  g09660(.a(n9267), .b(n3210), .O(n10608));
  andx  g09661(.a(n10209), .b(n10198), .O(n10609));
  orx   g09662(.a(n10209), .b(n10198), .O(n10610));
  andx  g09663(.a(n10610), .b(n10199), .O(n10611));
  orx   g09664(.a(n10611), .b(n10609), .O(n10612));
  andx  g09665(.a(n10612), .b(n10608), .O(n10613));
  invx  g09666(.a(n10608), .O(n10614));
  invx  g09667(.a(n10609), .O(n10615));
  andx  g09668(.a(n10204), .b(n10215), .O(n10616));
  orx   g09669(.a(n10616), .b(n10206), .O(n10617));
  andx  g09670(.a(n10617), .b(n10615), .O(n10618));
  andx  g09671(.a(n10618), .b(n10614), .O(n10619));
  orx   g09672(.a(n10619), .b(n10613), .O(n10620));
  orx   g09673(.a(n10620), .b(n10607), .O(n10621));
  orx   g09674(.a(n10605), .b(n10602), .O(n10622));
  orx   g09675(.a(n10598), .b(n10583), .O(n10623));
  andx  g09676(.a(n10623), .b(n10622), .O(n10624));
  orx   g09677(.a(n10618), .b(n10614), .O(n10625));
  orx   g09678(.a(n10612), .b(n10608), .O(n10626));
  andx  g09679(.a(n10626), .b(n10625), .O(n10627));
  orx   g09680(.a(n10627), .b(n10624), .O(n10628));
  andx  g09681(.a(n10628), .b(n10621), .O(n10629));
  andx  g09682(.a(n9470), .b(n3221), .O(n10630));
  invx  g09683(.a(n10630), .O(n10631));
  andx  g09684(.a(n10226), .b(n10237), .O(n10632));
  orx   g09685(.a(n10226), .b(n10237), .O(n10633));
  andx  g09686(.a(n10633), .b(n10221), .O(n10634));
  orx   g09687(.a(n10634), .b(n10632), .O(n10635));
  andx  g09688(.a(n10635), .b(n10631), .O(n10636));
  invx  g09689(.a(n10632), .O(n10637));
  andx  g09690(.a(n10231), .b(n10220), .O(n10638));
  orx   g09691(.a(n10638), .b(n10222), .O(n10639));
  andx  g09692(.a(n10639), .b(n10637), .O(n10640));
  andx  g09693(.a(n10640), .b(n10630), .O(n10641));
  orx   g09694(.a(n10641), .b(n10636), .O(n10642));
  andx  g09695(.a(n10642), .b(n10629), .O(n10643));
  andx  g09696(.a(n10627), .b(n10624), .O(n10644));
  andx  g09697(.a(n10620), .b(n10607), .O(n10645));
  orx   g09698(.a(n10645), .b(n10644), .O(n10646));
  orx   g09699(.a(n10640), .b(n10630), .O(n10647));
  orx   g09700(.a(n10635), .b(n10631), .O(n10648));
  andx  g09701(.a(n10648), .b(n10647), .O(n10649));
  andx  g09702(.a(n10649), .b(n10646), .O(n10650));
  orx   g09703(.a(n10650), .b(n10643), .O(n10651));
  andx  g09704(.a(n7902), .b(n3230), .O(n10652));
  andx  g09705(.a(n10253), .b(n10242), .O(n10653));
  invx  g09706(.a(n10653), .O(n10654));
  andx  g09707(.a(n10247), .b(n10259), .O(n10655));
  orx   g09708(.a(n10655), .b(n10249), .O(n10656));
  andx  g09709(.a(n10656), .b(n10654), .O(n10657));
  orx   g09710(.a(n10657), .b(n10652), .O(n10658));
  invx  g09711(.a(n10652), .O(n10659));
  orx   g09712(.a(n10253), .b(n10242), .O(n10660));
  andx  g09713(.a(n10660), .b(n10248), .O(n10661));
  orx   g09714(.a(n10661), .b(n10653), .O(n10662));
  orx   g09715(.a(n10662), .b(n10659), .O(n10663));
  andx  g09716(.a(n10663), .b(n10658), .O(n10664));
  orx   g09717(.a(n10664), .b(n10651), .O(n10665));
  orx   g09718(.a(n10649), .b(n10646), .O(n10666));
  orx   g09719(.a(n10642), .b(n10629), .O(n10667));
  andx  g09720(.a(n10667), .b(n10666), .O(n10668));
  andx  g09721(.a(n10662), .b(n10659), .O(n10669));
  andx  g09722(.a(n10657), .b(n10652), .O(n10670));
  orx   g09723(.a(n10670), .b(n10669), .O(n10671));
  orx   g09724(.a(n10671), .b(n10668), .O(n10672));
  andx  g09725(.a(n10672), .b(n10665), .O(n10673));
  andx  g09726(.a(n10356), .b(n3258), .O(n10674));
  invx  g09727(.a(n10674), .O(n10675));
  andx  g09728(.a(n10262), .b(n10259), .O(n10676));
  andx  g09729(.a(n10255), .b(n10242), .O(n10677));
  orx   g09730(.a(n10677), .b(n10676), .O(n10678));
  andx  g09731(.a(n10270), .b(n10678), .O(n10679));
  orx   g09732(.a(n10270), .b(n10678), .O(n10680));
  andx  g09733(.a(n10680), .b(n10265), .O(n10681));
  orx   g09734(.a(n10681), .b(n10679), .O(n10682));
  andx  g09735(.a(n10682), .b(n10675), .O(n10683));
  invx  g09736(.a(n10679), .O(n10684));
  andx  g09737(.a(n10275), .b(n10264), .O(n10685));
  orx   g09738(.a(n10685), .b(n10266), .O(n10686));
  andx  g09739(.a(n10686), .b(n10684), .O(n10687));
  andx  g09740(.a(n10687), .b(n10674), .O(n10688));
  orx   g09741(.a(n10688), .b(n10683), .O(n10689));
  andx  g09742(.a(n10689), .b(n10673), .O(n10690));
  invx  g09743(.a(n10690), .O(n10691));
  orx   g09744(.a(n10689), .b(n10673), .O(n10692));
  andx  g09745(.a(n10692), .b(n10691), .O(n10693));
  invx  g09746(.a(n10693), .O(n10694));
  andx  g09747(.a(n10323), .b(n10320), .O(n10695));
  orx   g09748(.a(n10695), .b(n10324), .O(n10696));
  invx  g09749(.a(n10696), .O(n10697));
  andx  g09750(.a(n826), .b(n4113), .O(n10703));
  invx  g09751(.a(n10703), .O(n10704));
  andx  g09752(.a(n10311), .b(n7676), .O(n10707));
  orx   g09753(.a(n10707), .b(n4113), .O(n10708));
  andx  g09754(.a(n10708), .b(n10314), .O(n10709));
  andx  g09755(.a(n10709), .b(n10704), .O(n10710));
  invx  g09756(.a(n10709), .O(n10711));
  andx  g09757(.a(n10711), .b(n10703), .O(n10712));
  orx   g09758(.a(n10712), .b(n10710), .O(n10713));
  invx  g09759(.a(n10713), .O(n10714));
  andx  g09760(.a(n2724), .b(n299), .O(n10715));
  invx  g09761(.a(n10715), .O(n10716));
  invx  g09762(.a(n10316), .O(n10717));
  andx  g09763(.a(n10717), .b(n10297), .O(n10718));
  orx   g09764(.a(n10718), .b(n602), .O(n10719));
  andx  g09765(.a(n10316), .b(n10298), .O(n10720));
  invx  g09766(.a(n10720), .O(n10721));
  andx  g09767(.a(n10721), .b(n10719), .O(n10722));
  invx  g09768(.a(n10722), .O(n10723));
  andx  g09769(.a(n10723), .b(n10716), .O(n10724));
  andx  g09770(.a(n10722), .b(n10715), .O(n10725));
  orx   g09771(.a(n10725), .b(n10724), .O(n10726));
  orx   g09772(.a(n10726), .b(n10714), .O(n10729));
  andx  g09773(.a(n10729), .b(n5793), .O(n10730));
  invx  g09774(.a(n10730), .O(n10731));
  andx  g09775(.a(n10731), .b(n10697), .O(n10732));
  andx  g09776(.a(n10730), .b(n10696), .O(n10733));
  orx   g09777(.a(n10733), .b(n10732), .O(n10734));
  andx  g09778(.a(n10734), .b(n10340), .O(n10735));
  invx  g09779(.a(n10735), .O(n10736));
  orx   g09780(.a(n10734), .b(n10340), .O(n10737));
  andx  g09781(.a(n10737), .b(n10736), .O(n10738));
  invx  g09782(.a(n10346), .O(n10739));
  andx  g09783(.a(n10345), .b(n10350), .O(n10740));
  orx   g09784(.a(n10740), .b(n10739), .O(n10741));
  andx  g09785(.a(n10741), .b(n10738), .O(n10742));
  invx  g09786(.a(n10742), .O(n10743));
  orx   g09787(.a(n10741), .b(n10738), .O(n10744));
  andx  g09788(.a(n10744), .b(n10743), .O(n10745));
  invx  g09789(.a(n10745), .O(n10746));
  andx  g09790(.a(n10352), .b(n10287), .O(n10747));
  invx  g09791(.a(n10747), .O(n10748));
  andx  g09792(.a(n10748), .b(n10746), .O(n10749));
  andx  g09793(.a(n10747), .b(n10745), .O(n10750));
  orx   g09794(.a(n10750), .b(n10749), .O(n10751));
  andx  g09795(.a(n10751), .b(n1790), .O(n10752));
  andx  g09796(.a(n10362), .b(n10367), .O(n10753));
  orx   g09797(.a(n10362), .b(n10367), .O(n10754));
  andx  g09798(.a(n10754), .b(n10357), .O(n10755));
  orx   g09799(.a(n10755), .b(n10753), .O(n10756));
  andx  g09800(.a(n10756), .b(n10752), .O(n10757));
  invx  g09801(.a(n10752), .O(n10758));
  invx  g09802(.a(n10753), .O(n10759));
  andx  g09803(.a(n10286), .b(n10281), .O(n10760));
  orx   g09804(.a(n10760), .b(n10358), .O(n10761));
  andx  g09805(.a(n10761), .b(n10759), .O(n10762));
  andx  g09806(.a(n10762), .b(n10758), .O(n10763));
  orx   g09807(.a(n10763), .b(n10757), .O(n10764));
  invx  g09808(.a(n10764), .O(n10765));
  orx   g09809(.a(n10765), .b(n10694), .O(n10766));
  orx   g09810(.a(n10764), .b(n10693), .O(n10767));
  andx  g09811(.a(n10767), .b(n10766), .O(po07));
  orx   g09812(.a(n10618), .b(n10624), .O(n10769));
  andx  g09813(.a(n10618), .b(n10624), .O(n10770));
  orx   g09814(.a(n10770), .b(n10614), .O(n10771));
  andx  g09815(.a(n10771), .b(n10769), .O(n10772));
  andx  g09816(.a(n9470), .b(n3210), .O(n10773));
  invx  g09817(.a(n10773), .O(n10774));
  andx  g09818(.a(n10774), .b(n10772), .O(n10775));
  andx  g09819(.a(n10612), .b(n10607), .O(n10776));
  orx   g09820(.a(n10612), .b(n10607), .O(n10777));
  andx  g09821(.a(n10777), .b(n10608), .O(n10778));
  orx   g09822(.a(n10778), .b(n10776), .O(n10779));
  andx  g09823(.a(n10779), .b(n9470), .O(n10780));
  orx   g09824(.a(n10780), .b(n10775), .O(n10781));
  andx  g09825(.a(n8852), .b(n3429), .O(n10782));
  invx  g09826(.a(n10782), .O(n10783));
  andx  g09827(.a(n10547), .b(n10544), .O(n10784));
  andx  g09828(.a(n10540), .b(n10527), .O(n10785));
  orx   g09829(.a(n10785), .b(n10784), .O(n10786));
  andx  g09830(.a(n10414), .b(n10786), .O(n10790));
  andx  g09831(.a(n10405), .b(n10407), .O(n10791));
  andx  g09832(.a(n10412), .b(n10400), .O(n10792));
  orx   g09833(.a(n10792), .b(n10791), .O(n10793));
  andx  g09834(.a(n10793), .b(n10549), .O(n10794));
  orx   g09835(.a(n10794), .b(n10790), .O(n10795));
  andx  g09836(.a(n10795), .b(n10560), .O(n10796));
  invx  g09837(.a(n10796), .O(n10797));
  orx   g09838(.a(n10793), .b(n10549), .O(n10798));
  orx   g09839(.a(n10414), .b(n10786), .O(n10799));
  andx  g09840(.a(n10799), .b(n10798), .O(n10800));
  orx   g09841(.a(n10800), .b(n10564), .O(n10801));
  orx   g09842(.a(n10564), .b(n10554), .O(n10802));
  andx  g09843(.a(n10802), .b(n10801), .O(n10803));
  andx  g09844(.a(n10803), .b(n10797), .O(n10804));
  orx   g09845(.a(n10804), .b(n10783), .O(n10805));
  andx  g09846(.a(n10795), .b(n10558), .O(n10806));
  andx  g09847(.a(n10558), .b(n10560), .O(n10807));
  orx   g09848(.a(n10807), .b(n10806), .O(n10808));
  orx   g09849(.a(n10808), .b(n10796), .O(n10809));
  orx   g09850(.a(n10809), .b(n10782), .O(n10810));
  andx  g09851(.a(n10810), .b(n10805), .O(n10811));
  andx  g09852(.a(n8603), .b(n3413), .O(n10812));
  andx  g09853(.a(n10528), .b(n10527), .O(n10813));
  andx  g09854(.a(n10538), .b(n10527), .O(n10814));
  andx  g09855(.a(n10538), .b(n10528), .O(n10815));
  orx   g09856(.a(n10815), .b(n10814), .O(n10816));
  orx   g09857(.a(n10816), .b(n10813), .O(n10817));
  andx  g09858(.a(n10817), .b(n10812), .O(n10818));
  orx   g09859(.a(n9680), .b(n4989), .O(n10819));
  invx  g09860(.a(n10813), .O(n10820));
  orx   g09861(.a(n10532), .b(n10544), .O(n10821));
  orx   g09862(.a(n10532), .b(n10534), .O(n10822));
  andx  g09863(.a(n10822), .b(n10821), .O(n10823));
  andx  g09864(.a(n10823), .b(n10820), .O(n10824));
  andx  g09865(.a(n10824), .b(n10819), .O(n10825));
  orx   g09866(.a(n10825), .b(n10818), .O(n10826));
  andx  g09867(.a(n8220), .b(n3721), .O(n10827));
  invx  g09868(.a(n10827), .O(n10828));
  andx  g09869(.a(n10474), .b(n10486), .O(n10829));
  andx  g09870(.a(n10473), .b(n10486), .O(n10830));
  orx   g09871(.a(n10830), .b(n10488), .O(n10831));
  orx   g09872(.a(n10831), .b(n10829), .O(n10832));
  andx  g09873(.a(n10832), .b(n10828), .O(n10833));
  invx  g09874(.a(n10829), .O(n10834));
  orx   g09875(.a(n10479), .b(n10466), .O(n10835));
  andx  g09876(.a(n10835), .b(n10481), .O(n10836));
  andx  g09877(.a(n10836), .b(n10834), .O(n10837));
  andx  g09878(.a(n10837), .b(n10827), .O(n10838));
  orx   g09879(.a(n10838), .b(n10833), .O(n10839));
  andx  g09880(.a(n7924), .b(n2724), .O(n10840));
  andx  g09881(.a(n2429), .b(n7982), .O(n10844));
  andx  g09882(.a(n10840), .b(n7931), .O(n10848));
  invx  g09883(.a(n10848), .O(n10849));
  andx  g09884(.a(n7959), .b(n8009), .O(n10850));
  orx   g09885(.a(n10850), .b(n10440), .O(n10851));
  andx  g09886(.a(n10851), .b(n10849), .O(n10852));
  invx  g09887(.a(n10844), .O(n10854));
  andx  g09888(.a(n8062), .b(n4114), .O(n10858));
  invx  g09889(.a(n10858), .O(n10859));
  andx  g09890(.a(n10433), .b(n10430), .O(n10860));
  orx   g09891(.a(n10433), .b(n10430), .O(n10861));
  andx  g09892(.a(n10861), .b(n7924), .O(n10862));
  orx   g09893(.a(n10862), .b(n10860), .O(n10863));
  andx  g09894(.a(n10863), .b(n10859), .O(n10864));
  invx  g09895(.a(n10864), .O(n10865));
  orx   g09896(.a(n10863), .b(n10859), .O(n10866));
  andx  g09897(.a(n10866), .b(n10865), .O(n10867));
  orx   g09898(.a(n10867), .b(n10844), .O(n10868));
  invx  g09899(.a(n10866), .O(n10869));
  orx   g09900(.a(n10869), .b(n10864), .O(n10870));
  orx   g09901(.a(n10870), .b(n10854), .O(n10871));
  andx  g09902(.a(n10871), .b(n10868), .O(n10872));
  andx  g09903(.a(n8131), .b(n4063), .O(n10873));
  invx  g09904(.a(n10873), .O(n10874));
  andx  g09905(.a(n10464), .b(n10421), .O(n10875));
  orx   g09906(.a(n10464), .b(n10421), .O(n10876));
  andx  g09907(.a(n10876), .b(n10415), .O(n10877));
  orx   g09908(.a(n10877), .b(n10875), .O(n10878));
  andx  g09909(.a(n10878), .b(n10874), .O(n10879));
  invx  g09910(.a(n10875), .O(n10880));
  andx  g09911(.a(n10457), .b(n10427), .O(n10881));
  orx   g09912(.a(n10881), .b(n10416), .O(n10882));
  andx  g09913(.a(n10882), .b(n10880), .O(n10883));
  andx  g09914(.a(n10883), .b(n10873), .O(n10884));
  orx   g09915(.a(n10884), .b(n10879), .O(n10885));
  andx  g09916(.a(n10885), .b(n10872), .O(n10886));
  andx  g09917(.a(n10870), .b(n10854), .O(n10887));
  andx  g09918(.a(n10867), .b(n10844), .O(n10888));
  orx   g09919(.a(n10888), .b(n10887), .O(n10889));
  orx   g09920(.a(n10883), .b(n10873), .O(n10890));
  orx   g09921(.a(n10878), .b(n10874), .O(n10891));
  andx  g09922(.a(n10891), .b(n10890), .O(n10892));
  andx  g09923(.a(n10892), .b(n10889), .O(n10893));
  orx   g09924(.a(n10893), .b(n10886), .O(n10894));
  andx  g09925(.a(n10894), .b(n10839), .O(n10895));
  orx   g09926(.a(n10837), .b(n10827), .O(n10896));
  orx   g09927(.a(n10832), .b(n10828), .O(n10897));
  andx  g09928(.a(n10897), .b(n10896), .O(n10898));
  orx   g09929(.a(n10892), .b(n10889), .O(n10899));
  orx   g09930(.a(n10885), .b(n10872), .O(n10900));
  andx  g09931(.a(n10900), .b(n10899), .O(n10901));
  andx  g09932(.a(n10901), .b(n10898), .O(n10902));
  orx   g09933(.a(n10902), .b(n10895), .O(n10903));
  andx  g09934(.a(n10515), .b(n10491), .O(n10904));
  orx   g09935(.a(n10515), .b(n10491), .O(n10905));
  andx  g09936(.a(n10905), .b(n10510), .O(n10906));
  orx   g09937(.a(n10906), .b(n10904), .O(n10907));
  andx  g09938(.a(n10907), .b(n8351), .O(n10908));
  invx  g09939(.a(n10904), .O(n10909));
  andx  g09940(.a(n10509), .b(n10522), .O(n10910));
  orx   g09941(.a(n10910), .b(n10516), .O(n10911));
  andx  g09942(.a(n10911), .b(n10909), .O(n10912));
  andx  g09943(.a(n8351), .b(n3645), .O(n10913));
  invx  g09944(.a(n10913), .O(n10914));
  andx  g09945(.a(n10914), .b(n10912), .O(n10915));
  orx   g09946(.a(n10915), .b(n10908), .O(n10916));
  andx  g09947(.a(n10916), .b(n10903), .O(n10917));
  orx   g09948(.a(n10901), .b(n10898), .O(n10918));
  orx   g09949(.a(n10894), .b(n10839), .O(n10919));
  andx  g09950(.a(n10919), .b(n10918), .O(n10920));
  orx   g09951(.a(n10912), .b(n9841), .O(n10921));
  orx   g09952(.a(n10913), .b(n10907), .O(n10922));
  andx  g09953(.a(n10922), .b(n10921), .O(n10923));
  andx  g09954(.a(n10923), .b(n10920), .O(n10924));
  orx   g09955(.a(n10924), .b(n10917), .O(n10925));
  orx   g09956(.a(n10925), .b(n10826), .O(n10926));
  orx   g09957(.a(n10824), .b(n10819), .O(n10927));
  orx   g09958(.a(n10817), .b(n10812), .O(n10928));
  andx  g09959(.a(n10928), .b(n10927), .O(n10929));
  orx   g09960(.a(n10923), .b(n10920), .O(n10930));
  orx   g09961(.a(n10916), .b(n10903), .O(n10931));
  andx  g09962(.a(n10931), .b(n10930), .O(n10932));
  orx   g09963(.a(n10932), .b(n10929), .O(n10933));
  andx  g09964(.a(n10933), .b(n10926), .O(n10934));
  orx   g09965(.a(n10549), .b(n10412), .O(n10935));
  andx  g09966(.a(n10549), .b(n10412), .O(n10936));
  orx   g09967(.a(n10936), .b(n10407), .O(n10937));
  andx  g09968(.a(n10937), .b(n10935), .O(n10938));
  orx   g09969(.a(n10938), .b(n10161), .O(n10939));
  andx  g09970(.a(n10786), .b(n10405), .O(n10940));
  orx   g09971(.a(n10786), .b(n10405), .O(n10941));
  andx  g09972(.a(n10941), .b(n10400), .O(n10942));
  orx   g09973(.a(n10942), .b(n10940), .O(n10943));
  andx  g09974(.a(n7907), .b(n3171), .O(n10944));
  orx   g09975(.a(n10944), .b(n10943), .O(n10945));
  andx  g09976(.a(n10945), .b(n10939), .O(n10946));
  orx   g09977(.a(n10946), .b(n10934), .O(n10947));
  andx  g09978(.a(n10932), .b(n10929), .O(n10948));
  andx  g09979(.a(n10925), .b(n10826), .O(n10949));
  orx   g09980(.a(n10949), .b(n10948), .O(n10950));
  andx  g09981(.a(n10943), .b(n7907), .O(n10951));
  orx   g09982(.a(n10161), .b(n3418), .O(n10952));
  andx  g09983(.a(n10952), .b(n10938), .O(n10953));
  orx   g09984(.a(n10953), .b(n10951), .O(n10954));
  orx   g09985(.a(n10954), .b(n10950), .O(n10955));
  andx  g09986(.a(n10955), .b(n10947), .O(n10956));
  andx  g09987(.a(n10956), .b(n10811), .O(n10957));
  andx  g09988(.a(n10809), .b(n10782), .O(n10958));
  andx  g09989(.a(n10804), .b(n10783), .O(n10959));
  orx   g09990(.a(n10959), .b(n10958), .O(n10960));
  andx  g09991(.a(n10954), .b(n10950), .O(n10961));
  andx  g09992(.a(n10946), .b(n10934), .O(n10962));
  orx   g09993(.a(n10962), .b(n10961), .O(n10963));
  andx  g09994(.a(n10963), .b(n10960), .O(n10964));
  orx   g09995(.a(n10964), .b(n10957), .O(n10965));
  andx  g09996(.a(n10574), .b(n10397), .O(n10966));
  orx   g09997(.a(n10574), .b(n10397), .O(n10967));
  andx  g09998(.a(n10967), .b(n10370), .O(n10968));
  orx   g09999(.a(n10968), .b(n10966), .O(n10969));
  andx  g10000(.a(n10969), .b(n9050), .O(n10970));
  orx   g10001(.a(n10581), .b(n10392), .O(n10971));
  andx  g10002(.a(n10581), .b(n10392), .O(n10972));
  orx   g10003(.a(n10972), .b(n10371), .O(n10973));
  andx  g10004(.a(n10973), .b(n10971), .O(n10974));
  orx   g10005(.a(n10585), .b(n3183), .O(n10975));
  andx  g10006(.a(n10975), .b(n10974), .O(n10976));
  orx   g10007(.a(n10976), .b(n10970), .O(n10977));
  andx  g10008(.a(n10977), .b(n10965), .O(n10978));
  orx   g10009(.a(n10963), .b(n10960), .O(n10979));
  orx   g10010(.a(n10956), .b(n10811), .O(n10980));
  andx  g10011(.a(n10980), .b(n10979), .O(n10981));
  orx   g10012(.a(n10974), .b(n10585), .O(n10982));
  andx  g10013(.a(n9050), .b(n3180), .O(n10983));
  orx   g10014(.a(n10983), .b(n10969), .O(n10984));
  andx  g10015(.a(n10984), .b(n10982), .O(n10985));
  andx  g10016(.a(n10985), .b(n10981), .O(n10986));
  orx   g10017(.a(n10986), .b(n10978), .O(n10987));
  andx  g10018(.a(n9267), .b(n3284), .O(n10988));
  invx  g10019(.a(n10988), .O(n10989));
  andx  g10020(.a(n10590), .b(n10602), .O(n10990));
  invx  g10021(.a(n10990), .O(n10991));
  andx  g10022(.a(n10596), .b(n10583), .O(n10992));
  orx   g10023(.a(n10992), .b(n10586), .O(n10993));
  andx  g10024(.a(n10993), .b(n10991), .O(n10994));
  orx   g10025(.a(n10994), .b(n10989), .O(n10995));
  orx   g10026(.a(n10590), .b(n10602), .O(n10996));
  andx  g10027(.a(n10996), .b(n10592), .O(n10997));
  orx   g10028(.a(n10997), .b(n10990), .O(n10998));
  orx   g10029(.a(n10998), .b(n10988), .O(n10999));
  andx  g10030(.a(n10999), .b(n10995), .O(n11000));
  andx  g10031(.a(n11000), .b(n10987), .O(n11001));
  orx   g10032(.a(n10985), .b(n10981), .O(n11002));
  orx   g10033(.a(n10977), .b(n10965), .O(n11003));
  andx  g10034(.a(n11003), .b(n11002), .O(n11004));
  andx  g10035(.a(n10998), .b(n10988), .O(n11005));
  andx  g10036(.a(n10994), .b(n10989), .O(n11006));
  orx   g10037(.a(n11006), .b(n11005), .O(n11007));
  andx  g10038(.a(n11007), .b(n11004), .O(n11008));
  orx   g10039(.a(n11008), .b(n11001), .O(n11009));
  andx  g10040(.a(n11009), .b(n10781), .O(n11010));
  orx   g10041(.a(n10773), .b(n10779), .O(n11011));
  invx  g10042(.a(n9470), .O(n11012));
  orx   g10043(.a(n10772), .b(n11012), .O(n11013));
  andx  g10044(.a(n11013), .b(n11011), .O(n11014));
  orx   g10045(.a(n11007), .b(n11004), .O(n11015));
  orx   g10046(.a(n11000), .b(n10987), .O(n11016));
  andx  g10047(.a(n11016), .b(n11015), .O(n11017));
  andx  g10048(.a(n11017), .b(n11014), .O(n11018));
  orx   g10049(.a(n11018), .b(n11010), .O(n11019));
  andx  g10050(.a(n10635), .b(n10646), .O(n11020));
  invx  g10051(.a(n11020), .O(n11021));
  andx  g10052(.a(n10640), .b(n10629), .O(n11022));
  orx   g10053(.a(n11022), .b(n10631), .O(n11023));
  andx  g10054(.a(n11023), .b(n11021), .O(n11024));
  andx  g10055(.a(n7902), .b(n3221), .O(n11025));
  invx  g10056(.a(n11025), .O(n11026));
  andx  g10057(.a(n11026), .b(n11024), .O(n11027));
  orx   g10058(.a(n10635), .b(n10646), .O(n11028));
  andx  g10059(.a(n11028), .b(n10630), .O(n11029));
  orx   g10060(.a(n11029), .b(n11020), .O(n11030));
  andx  g10061(.a(n11025), .b(n11030), .O(n11031));
  orx   g10062(.a(n11031), .b(n11027), .O(n11032));
  orx   g10063(.a(n11032), .b(n11019), .O(n11033));
  andx  g10064(.a(n11032), .b(n11019), .O(n11034));
  invx  g10065(.a(n11034), .O(n11035));
  andx  g10066(.a(n11035), .b(n11033), .O(n11036));
  andx  g10067(.a(n10662), .b(n10651), .O(n11037));
  orx   g10068(.a(n10662), .b(n10651), .O(n11038));
  andx  g10069(.a(n11038), .b(n10652), .O(n11039));
  orx   g10070(.a(n11039), .b(n11037), .O(n11040));
  andx  g10071(.a(n11040), .b(n10356), .O(n11041));
  invx  g10072(.a(n11037), .O(n11042));
  andx  g10073(.a(n10657), .b(n10668), .O(n11043));
  orx   g10074(.a(n11043), .b(n10659), .O(n11044));
  andx  g10075(.a(n11044), .b(n11042), .O(n11045));
  andx  g10076(.a(n10356), .b(n3230), .O(n11046));
  invx  g10077(.a(n11046), .O(n11047));
  andx  g10078(.a(n11047), .b(n11045), .O(n11048));
  orx   g10079(.a(n11048), .b(n11041), .O(n11049));
  andx  g10080(.a(n11049), .b(n11036), .O(n11050));
  invx  g10081(.a(n11033), .O(n11051));
  orx   g10082(.a(n11034), .b(n11051), .O(n11052));
  invx  g10083(.a(n10356), .O(n11053));
  orx   g10084(.a(n11045), .b(n11053), .O(n11054));
  orx   g10085(.a(n11046), .b(n11040), .O(n11055));
  andx  g10086(.a(n11055), .b(n11054), .O(n11056));
  andx  g10087(.a(n11056), .b(n11052), .O(n11057));
  orx   g10088(.a(n11057), .b(n11050), .O(n11058));
  andx  g10089(.a(n10671), .b(n10668), .O(n11059));
  andx  g10090(.a(n10664), .b(n10651), .O(n11060));
  orx   g10091(.a(n11060), .b(n11059), .O(n11061));
  andx  g10092(.a(n10682), .b(n11061), .O(n11062));
  invx  g10093(.a(n11062), .O(n11063));
  andx  g10094(.a(n10687), .b(n10673), .O(n11064));
  orx   g10095(.a(n11064), .b(n10675), .O(n11065));
  andx  g10096(.a(n11065), .b(n11063), .O(n11066));
  andx  g10097(.a(n10751), .b(n3258), .O(n11067));
  invx  g10098(.a(n11067), .O(n11068));
  andx  g10099(.a(n11068), .b(n11066), .O(n11069));
  orx   g10100(.a(n10682), .b(n11061), .O(n11070));
  andx  g10101(.a(n11070), .b(n10674), .O(n11071));
  orx   g10102(.a(n11071), .b(n11062), .O(n11072));
  andx  g10103(.a(n11067), .b(n11072), .O(n11073));
  orx   g10104(.a(n11073), .b(n11069), .O(n11074));
  invx  g10105(.a(n11074), .O(n11075));
  andx  g10106(.a(n11075), .b(n11058), .O(n11076));
  orx   g10107(.a(n11056), .b(n11052), .O(n11077));
  orx   g10108(.a(n11049), .b(n11036), .O(n11078));
  andx  g10109(.a(n11078), .b(n11077), .O(n11079));
  andx  g10110(.a(n11074), .b(n11079), .O(n11080));
  orx   g10111(.a(n11080), .b(n11076), .O(n11081));
  andx  g10112(.a(n10747), .b(n10746), .O(n11082));
  invx  g10113(.a(n11082), .O(n11083));
  andx  g10114(.a(n10723), .b(n10713), .O(n11084));
  andx  g10115(.a(n10715), .b(n10713), .O(n11085));
  andx  g10116(.a(n10723), .b(n10715), .O(n11086));
  orx   g10117(.a(n11086), .b(n11085), .O(n11087));
  orx   g10118(.a(n11087), .b(n11084), .O(n11088));
  andx  g10119(.a(n10709), .b(n10303), .O(n11093));
  orx   g10120(.a(n11093), .b(n5878), .O(n11094));
  andx  g10121(.a(n10711), .b(n4114), .O(n11095));
  invx  g10122(.a(n11095), .O(n11096));
  andx  g10123(.a(n11096), .b(n11094), .O(n11097));
  invx  g10124(.a(n11097), .O(n11098));
  andx  g10125(.a(n11098), .b(n2429), .O(n11099));
  invx  g10126(.a(n11099), .O(n11100));
  andx  g10127(.a(n2429), .b(n11100), .O(n11102));
  invx  g10128(.a(n11102), .O(n11103));
  andx  g10129(.a(n11103), .b(n11088), .O(n11104));
  invx  g10130(.a(n11088), .O(n11105));
  andx  g10131(.a(n11102), .b(n11105), .O(n11106));
  orx   g10132(.a(n11106), .b(n11104), .O(n11107));
  invx  g10133(.a(n11107), .O(n11108));
  andx  g10134(.a(n10731), .b(n10696), .O(n11109));
  orx   g10135(.a(n11109), .b(n10735), .O(n11110));
  andx  g10136(.a(n10741), .b(n10737), .O(n11111));
  orx   g10137(.a(n11111), .b(n11110), .O(n11112));
  andx  g10138(.a(n11112), .b(n11108), .O(n11113));
  invx  g10139(.a(n11113), .O(n11114));
  orx   g10140(.a(n11112), .b(n11108), .O(n11115));
  andx  g10141(.a(n11115), .b(n11114), .O(n11116));
  andx  g10142(.a(n11116), .b(n11083), .O(n11117));
  invx  g10143(.a(n11116), .O(n11118));
  andx  g10144(.a(n11118), .b(n11082), .O(n11119));
  orx   g10145(.a(n11119), .b(n11117), .O(n11120));
  andx  g10146(.a(n10756), .b(n10694), .O(n11121));
  orx   g10147(.a(n10756), .b(n10694), .O(n11122));
  andx  g10148(.a(n11122), .b(n10752), .O(n11123));
  orx   g10149(.a(n11123), .b(n11121), .O(n11124));
  andx  g10150(.a(n11124), .b(n11120), .O(n11125));
  invx  g10151(.a(n11125), .O(n11126));
  andx  g10152(.a(n11120), .b(n1790), .O(n11127));
  orx   g10153(.a(n11127), .b(n11124), .O(n11128));
  andx  g10154(.a(n11128), .b(n11126), .O(n11129));
  orx   g10155(.a(n11129), .b(n11081), .O(n11130));
  invx  g10156(.a(n11081), .O(n11131));
  invx  g10157(.a(n11129), .O(n11132));
  orx   g10158(.a(n11132), .b(n11131), .O(n11133));
  andx  g10159(.a(n11133), .b(n11130), .O(po08));
  andx  g10160(.a(n8351), .b(n3721), .O(n11135));
  andx  g10161(.a(n10894), .b(n10832), .O(n11136));
  invx  g10162(.a(n11136), .O(n11137));
  andx  g10163(.a(n10901), .b(n10837), .O(n11138));
  orx   g10164(.a(n11138), .b(n10828), .O(n11139));
  andx  g10165(.a(n11139), .b(n11137), .O(n11140));
  orx   g10166(.a(n11140), .b(n11135), .O(n11141));
  invx  g10167(.a(n11135), .O(n11142));
  orx   g10168(.a(n10894), .b(n10832), .O(n11143));
  andx  g10169(.a(n11143), .b(n10827), .O(n11144));
  orx   g10170(.a(n11144), .b(n11136), .O(n11145));
  orx   g10171(.a(n11145), .b(n11142), .O(n11146));
  andx  g10172(.a(n11146), .b(n11141), .O(n11147));
  andx  g10173(.a(n2429), .b(n8062), .O(n11150));
  orx   g10174(.a(n7624), .b(n11150), .O(n11154));
  invx  g10175(.a(n10852), .O(n11155));
  andx  g10176(.a(n11155), .b(n10840), .O(n11156));
  andx  g10177(.a(n2724), .b(n4490), .O(n11157));
  andx  g10178(.a(n11157), .b(n7924), .O(n11158));
  orx   g10179(.a(n11158), .b(n11155), .O(n11159));
  andx  g10180(.a(n11159), .b(n7982), .O(n11160));
  orx   g10181(.a(n11160), .b(n11156), .O(n11161));
  invx  g10182(.a(n11154), .O(n11164));
  andx  g10183(.a(n8131), .b(n4114), .O(n11168));
  invx  g10184(.a(n11168), .O(n11169));
  andx  g10185(.a(n10863), .b(n10844), .O(n11170));
  orx   g10186(.a(n10863), .b(n10844), .O(n11171));
  andx  g10187(.a(n11171), .b(n10858), .O(n11172));
  orx   g10188(.a(n11172), .b(n11170), .O(n11173));
  andx  g10189(.a(n11173), .b(n11169), .O(n11174));
  invx  g10190(.a(n11174), .O(n11175));
  orx   g10191(.a(n11173), .b(n11169), .O(n11176));
  andx  g10192(.a(n11176), .b(n11175), .O(n11177));
  orx   g10193(.a(n11177), .b(n11154), .O(n11178));
  invx  g10194(.a(n11176), .O(n11179));
  orx   g10195(.a(n11179), .b(n11174), .O(n11180));
  orx   g10196(.a(n11180), .b(n11164), .O(n11181));
  andx  g10197(.a(n11181), .b(n11178), .O(n11182));
  andx  g10198(.a(n10878), .b(n10889), .O(n11183));
  orx   g10199(.a(n10878), .b(n10889), .O(n11184));
  andx  g10200(.a(n11184), .b(n10873), .O(n11185));
  orx   g10201(.a(n11185), .b(n11183), .O(n11186));
  andx  g10202(.a(n11186), .b(n8220), .O(n11187));
  invx  g10203(.a(n11183), .O(n11188));
  andx  g10204(.a(n10883), .b(n10872), .O(n11189));
  orx   g10205(.a(n11189), .b(n10874), .O(n11190));
  andx  g10206(.a(n11190), .b(n11188), .O(n11191));
  andx  g10207(.a(n8220), .b(n4063), .O(n11192));
  invx  g10208(.a(n11192), .O(n11193));
  andx  g10209(.a(n11193), .b(n11191), .O(n11194));
  orx   g10210(.a(n11194), .b(n11187), .O(n11195));
  andx  g10211(.a(n11195), .b(n11182), .O(n11196));
  andx  g10212(.a(n11180), .b(n11164), .O(n11197));
  andx  g10213(.a(n11177), .b(n11154), .O(n11198));
  orx   g10214(.a(n11198), .b(n11197), .O(n11199));
  orx   g10215(.a(n11191), .b(n8675), .O(n11200));
  orx   g10216(.a(n11192), .b(n11186), .O(n11201));
  andx  g10217(.a(n11201), .b(n11200), .O(n11202));
  andx  g10218(.a(n11202), .b(n11199), .O(n11203));
  orx   g10219(.a(n11203), .b(n11196), .O(n11204));
  orx   g10220(.a(n11204), .b(n11147), .O(n11205));
  andx  g10221(.a(n11145), .b(n11142), .O(n11206));
  andx  g10222(.a(n11140), .b(n11135), .O(n11207));
  orx   g10223(.a(n11207), .b(n11206), .O(n11208));
  orx   g10224(.a(n11202), .b(n11199), .O(n11209));
  orx   g10225(.a(n11195), .b(n11182), .O(n11210));
  andx  g10226(.a(n11210), .b(n11209), .O(n11211));
  orx   g10227(.a(n11211), .b(n11208), .O(n11212));
  andx  g10228(.a(n11212), .b(n11205), .O(n11213));
  orx   g10229(.a(n10915), .b(n10903), .O(n11214));
  andx  g10230(.a(n11214), .b(n10921), .O(n11215));
  orx   g10231(.a(n11215), .b(n9680), .O(n11216));
  andx  g10232(.a(n10922), .b(n10920), .O(n11217));
  orx   g10233(.a(n11217), .b(n10908), .O(n11218));
  andx  g10234(.a(n8603), .b(n3645), .O(n11219));
  orx   g10235(.a(n11219), .b(n11218), .O(n11220));
  andx  g10236(.a(n11220), .b(n11216), .O(n11221));
  orx   g10237(.a(n11221), .b(n11213), .O(n11222));
  andx  g10238(.a(n11211), .b(n11208), .O(n11223));
  andx  g10239(.a(n11204), .b(n11147), .O(n11224));
  orx   g10240(.a(n11224), .b(n11223), .O(n11225));
  andx  g10241(.a(n11218), .b(n8603), .O(n11226));
  invx  g10242(.a(n11219), .O(n11227));
  andx  g10243(.a(n11227), .b(n11215), .O(n11228));
  orx   g10244(.a(n11228), .b(n11226), .O(n11229));
  orx   g10245(.a(n11229), .b(n11225), .O(n11230));
  andx  g10246(.a(n11230), .b(n11222), .O(n11231));
  andx  g10247(.a(n7907), .b(n3413), .O(n11232));
  andx  g10248(.a(n10932), .b(n10817), .O(n11233));
  orx   g10249(.a(n10932), .b(n10817), .O(n11234));
  andx  g10250(.a(n11234), .b(n10812), .O(n11235));
  orx   g10251(.a(n11235), .b(n11233), .O(n11236));
  andx  g10252(.a(n11236), .b(n11232), .O(n11237));
  invx  g10253(.a(n11232), .O(n11238));
  invx  g10254(.a(n11233), .O(n11239));
  andx  g10255(.a(n10925), .b(n10824), .O(n11240));
  orx   g10256(.a(n11240), .b(n10819), .O(n11241));
  andx  g10257(.a(n11241), .b(n11239), .O(n11242));
  andx  g10258(.a(n11242), .b(n11238), .O(n11243));
  orx   g10259(.a(n11243), .b(n11237), .O(n11244));
  orx   g10260(.a(n11244), .b(n11231), .O(n11245));
  andx  g10261(.a(n11229), .b(n11225), .O(n11246));
  andx  g10262(.a(n11221), .b(n11213), .O(n11247));
  orx   g10263(.a(n11247), .b(n11246), .O(n11248));
  orx   g10264(.a(n11242), .b(n11238), .O(n11249));
  orx   g10265(.a(n11236), .b(n11232), .O(n11250));
  andx  g10266(.a(n11250), .b(n11249), .O(n11251));
  orx   g10267(.a(n11251), .b(n11248), .O(n11252));
  andx  g10268(.a(n11252), .b(n11245), .O(n11253));
  andx  g10269(.a(n10945), .b(n10934), .O(n11254));
  orx   g10270(.a(n11254), .b(n10951), .O(n11255));
  andx  g10271(.a(n11255), .b(n8852), .O(n11256));
  orx   g10272(.a(n10953), .b(n10950), .O(n11257));
  andx  g10273(.a(n11257), .b(n10939), .O(n11258));
  andx  g10274(.a(n8849), .b(n8843), .O(n11259));
  orx   g10275(.a(n11259), .b(n7880), .O(n11260));
  orx   g10276(.a(n11260), .b(n3418), .O(n11261));
  andx  g10277(.a(n11261), .b(n11258), .O(n11262));
  orx   g10278(.a(n11262), .b(n11256), .O(n11263));
  andx  g10279(.a(n11263), .b(n11253), .O(n11264));
  andx  g10280(.a(n11251), .b(n11248), .O(n11265));
  andx  g10281(.a(n11244), .b(n11231), .O(n11266));
  orx   g10282(.a(n11266), .b(n11265), .O(n11267));
  orx   g10283(.a(n11258), .b(n11260), .O(n11268));
  andx  g10284(.a(n8852), .b(n3171), .O(n11269));
  orx   g10285(.a(n11269), .b(n11255), .O(n11270));
  andx  g10286(.a(n11270), .b(n11268), .O(n11271));
  andx  g10287(.a(n11271), .b(n11267), .O(n11272));
  orx   g10288(.a(n11272), .b(n11264), .O(n11273));
  orx   g10289(.a(n10585), .b(n3297), .O(n11274));
  andx  g10290(.a(n10956), .b(n10809), .O(n11275));
  orx   g10291(.a(n10956), .b(n10809), .O(n11276));
  andx  g10292(.a(n11276), .b(n10782), .O(n11277));
  orx   g10293(.a(n11277), .b(n11275), .O(n11278));
  andx  g10294(.a(n11278), .b(n11274), .O(n11279));
  andx  g10295(.a(n9050), .b(n3429), .O(n11280));
  orx   g10296(.a(n10963), .b(n10804), .O(n11281));
  andx  g10297(.a(n10963), .b(n10804), .O(n11282));
  orx   g10298(.a(n11282), .b(n10783), .O(n11283));
  andx  g10299(.a(n11283), .b(n11281), .O(n11284));
  andx  g10300(.a(n11284), .b(n11280), .O(n11285));
  orx   g10301(.a(n11285), .b(n11279), .O(n11286));
  andx  g10302(.a(n11286), .b(n11273), .O(n11287));
  orx   g10303(.a(n11271), .b(n11267), .O(n11288));
  orx   g10304(.a(n11263), .b(n11253), .O(n11289));
  andx  g10305(.a(n11289), .b(n11288), .O(n11290));
  orx   g10306(.a(n11284), .b(n11280), .O(n11291));
  orx   g10307(.a(n11278), .b(n11274), .O(n11292));
  andx  g10308(.a(n11292), .b(n11291), .O(n11293));
  andx  g10309(.a(n11293), .b(n11290), .O(n11294));
  orx   g10310(.a(n11294), .b(n11287), .O(n11295));
  orx   g10311(.a(n10976), .b(n10965), .O(n11296));
  andx  g10312(.a(n11296), .b(n10982), .O(n11297));
  orx   g10313(.a(n11297), .b(n9266), .O(n11298));
  andx  g10314(.a(n10984), .b(n10981), .O(n11299));
  orx   g10315(.a(n11299), .b(n10970), .O(n11300));
  orx   g10316(.a(n9266), .b(n3183), .O(n11301));
  invx  g10317(.a(n11301), .O(n11302));
  orx   g10318(.a(n11302), .b(n11300), .O(n11303));
  andx  g10319(.a(n11303), .b(n11298), .O(n11304));
  orx   g10320(.a(n11304), .b(n11295), .O(n11305));
  orx   g10321(.a(n11293), .b(n11290), .O(n11306));
  orx   g10322(.a(n11286), .b(n11273), .O(n11307));
  andx  g10323(.a(n11307), .b(n11306), .O(n11308));
  andx  g10324(.a(n11300), .b(n9267), .O(n11309));
  andx  g10325(.a(n11301), .b(n11297), .O(n11310));
  orx   g10326(.a(n11310), .b(n11309), .O(n11311));
  orx   g10327(.a(n11311), .b(n11308), .O(n11312));
  andx  g10328(.a(n11312), .b(n11305), .O(n11313));
  andx  g10329(.a(n9470), .b(n3284), .O(n11314));
  andx  g10330(.a(n10998), .b(n11004), .O(n11315));
  orx   g10331(.a(n10998), .b(n11004), .O(n11316));
  andx  g10332(.a(n11316), .b(n10988), .O(n11317));
  orx   g10333(.a(n11317), .b(n11315), .O(n11318));
  andx  g10334(.a(n11318), .b(n11314), .O(n11319));
  invx  g10335(.a(n11314), .O(n11320));
  orx   g10336(.a(n10994), .b(n10987), .O(n11321));
  andx  g10337(.a(n10994), .b(n10987), .O(n11322));
  orx   g10338(.a(n11322), .b(n10989), .O(n11323));
  andx  g10339(.a(n11323), .b(n11321), .O(n11324));
  andx  g10340(.a(n11324), .b(n11320), .O(n11325));
  orx   g10341(.a(n11325), .b(n11319), .O(n11326));
  orx   g10342(.a(n11326), .b(n11313), .O(n11327));
  andx  g10343(.a(n11311), .b(n11308), .O(n11328));
  andx  g10344(.a(n11304), .b(n11295), .O(n11329));
  orx   g10345(.a(n11329), .b(n11328), .O(n11330));
  orx   g10346(.a(n11324), .b(n11320), .O(n11331));
  orx   g10347(.a(n11318), .b(n11314), .O(n11332));
  andx  g10348(.a(n11332), .b(n11331), .O(n11333));
  orx   g10349(.a(n11333), .b(n11330), .O(n11334));
  andx  g10350(.a(n11334), .b(n11327), .O(n11335));
  andx  g10351(.a(n11009), .b(n11011), .O(n11336));
  orx   g10352(.a(n11336), .b(n10780), .O(n11337));
  andx  g10353(.a(n11337), .b(n7902), .O(n11338));
  orx   g10354(.a(n11017), .b(n10775), .O(n11339));
  andx  g10355(.a(n11339), .b(n11013), .O(n11340));
  andx  g10356(.a(n7902), .b(n3210), .O(n11341));
  invx  g10357(.a(n11341), .O(n11342));
  andx  g10358(.a(n11342), .b(n11340), .O(n11343));
  orx   g10359(.a(n11343), .b(n11338), .O(n11344));
  andx  g10360(.a(n11344), .b(n11335), .O(n11345));
  andx  g10361(.a(n11333), .b(n11330), .O(n11346));
  andx  g10362(.a(n11326), .b(n11313), .O(n11347));
  orx   g10363(.a(n11347), .b(n11346), .O(n11348));
  invx  g10364(.a(n7902), .O(n11349));
  orx   g10365(.a(n11340), .b(n11349), .O(n11350));
  orx   g10366(.a(n11341), .b(n11337), .O(n11351));
  andx  g10367(.a(n11351), .b(n11350), .O(n11352));
  andx  g10368(.a(n11352), .b(n11348), .O(n11353));
  orx   g10369(.a(n11353), .b(n11345), .O(n11354));
  andx  g10370(.a(n11030), .b(n11019), .O(n11355));
  orx   g10371(.a(n11030), .b(n11019), .O(n11356));
  andx  g10372(.a(n11356), .b(n11025), .O(n11357));
  orx   g10373(.a(n11357), .b(n11355), .O(n11358));
  andx  g10374(.a(n10356), .b(n3221), .O(n11359));
  orx   g10375(.a(n11359), .b(n11358), .O(n11360));
  orx   g10376(.a(n11017), .b(n11014), .O(n11361));
  orx   g10377(.a(n11009), .b(n10781), .O(n11362));
  andx  g10378(.a(n11362), .b(n11361), .O(n11363));
  orx   g10379(.a(n11024), .b(n11363), .O(n11364));
  andx  g10380(.a(n11024), .b(n11363), .O(n11365));
  orx   g10381(.a(n11365), .b(n11026), .O(n11366));
  andx  g10382(.a(n11366), .b(n11364), .O(n11367));
  invx  g10383(.a(n11359), .O(n11368));
  orx   g10384(.a(n11368), .b(n11367), .O(n11369));
  andx  g10385(.a(n11369), .b(n11360), .O(n11370));
  andx  g10386(.a(n11370), .b(n11354), .O(n11371));
  orx   g10387(.a(n11352), .b(n11348), .O(n11372));
  orx   g10388(.a(n11344), .b(n11335), .O(n11373));
  andx  g10389(.a(n11373), .b(n11372), .O(n11374));
  andx  g10390(.a(n11368), .b(n11367), .O(n11375));
  andx  g10391(.a(n11359), .b(n11358), .O(n11376));
  orx   g10392(.a(n11376), .b(n11375), .O(n11377));
  andx  g10393(.a(n11377), .b(n11374), .O(n11378));
  orx   g10394(.a(n11378), .b(n11371), .O(n11379));
  invx  g10395(.a(n10751), .O(n11380));
  orx   g10396(.a(n11048), .b(n11036), .O(n11381));
  andx  g10397(.a(n11381), .b(n11054), .O(n11382));
  orx   g10398(.a(n11382), .b(n11380), .O(n11383));
  andx  g10399(.a(n11055), .b(n11052), .O(n11384));
  orx   g10400(.a(n11384), .b(n11041), .O(n11385));
  andx  g10401(.a(n10751), .b(n3230), .O(n11386));
  orx   g10402(.a(n11386), .b(n11385), .O(n11387));
  andx  g10403(.a(n11387), .b(n11383), .O(n11388));
  orx   g10404(.a(n11388), .b(n11379), .O(n11389));
  orx   g10405(.a(n11377), .b(n11374), .O(n11390));
  orx   g10406(.a(n11370), .b(n11354), .O(n11391));
  andx  g10407(.a(n11391), .b(n11390), .O(n11392));
  andx  g10408(.a(n11385), .b(n10751), .O(n11393));
  invx  g10409(.a(n11386), .O(n11394));
  andx  g10410(.a(n11394), .b(n11382), .O(n11395));
  orx   g10411(.a(n11395), .b(n11393), .O(n11396));
  orx   g10412(.a(n11396), .b(n11392), .O(n11397));
  andx  g10413(.a(n11397), .b(n11389), .O(n11398));
  andx  g10414(.a(n11072), .b(n11079), .O(n11399));
  invx  g10415(.a(n11399), .O(n11400));
  andx  g10416(.a(n11066), .b(n11058), .O(n11401));
  orx   g10417(.a(n11401), .b(n11068), .O(n11402));
  andx  g10418(.a(n11402), .b(n11400), .O(n11403));
  andx  g10419(.a(n11120), .b(n3258), .O(n11404));
  invx  g10420(.a(n11404), .O(n11405));
  andx  g10421(.a(n11405), .b(n11403), .O(n11406));
  orx   g10422(.a(n11072), .b(n11079), .O(n11407));
  andx  g10423(.a(n11407), .b(n11067), .O(n11408));
  orx   g10424(.a(n11408), .b(n11399), .O(n11409));
  andx  g10425(.a(n11404), .b(n11409), .O(n11410));
  orx   g10426(.a(n11410), .b(n11406), .O(n11411));
  orx   g10427(.a(n11411), .b(n11398), .O(n11412));
  andx  g10428(.a(n11411), .b(n11398), .O(n11413));
  invx  g10429(.a(n11413), .O(n11414));
  andx  g10430(.a(n11414), .b(n11412), .O(n11415));
  invx  g10431(.a(n11415), .O(n11416));
  andx  g10432(.a(n11102), .b(n11088), .O(n11417));
  invx  g10433(.a(n11417), .O(n11418));
  andx  g10434(.a(n11418), .b(n2723), .O(n11419));
  andx  g10435(.a(n11417), .b(n2724), .O(n11420));
  orx   g10436(.a(n11420), .b(n11419), .O(n11421));
  orx   g10437(.a(n82), .b(n11097), .O(n11423));
  andx  g10438(.a(n11157), .b(n827), .O(n11424));
  invx  g10439(.a(n11424), .O(n11425));
  andx  g10440(.a(n11425), .b(n11423), .O(n11426));
  andx  g10441(.a(n10345), .b(n7658), .O(n11427));
  andx  g10442(.a(n11427), .b(n7724), .O(n11428));
  orx   g10443(.a(n11428), .b(n10739), .O(n11429));
  andx  g10444(.a(n11429), .b(n10737), .O(n11430));
  orx   g10445(.a(n11430), .b(n11110), .O(n11431));
  andx  g10446(.a(n11431), .b(n11107), .O(n11432));
  andx  g10447(.a(n11107), .b(n10737), .O(n11433));
  andx  g10448(.a(n10345), .b(n7724), .O(n11434));
  andx  g10449(.a(n11434), .b(n11433), .O(n11435));
  andx  g10450(.a(n11435), .b(n7656), .O(n11436));
  orx   g10451(.a(n11436), .b(n11432), .O(n11437));
  andx  g10452(.a(n11116), .b(n11082), .O(n11438));
  invx  g10453(.a(n11438), .O(n11439));
  andx  g10454(.a(n11439), .b(n11437), .O(n11440));
  invx  g10455(.a(n11440), .O(n11441));
  orx   g10456(.a(n11439), .b(n11437), .O(n11442));
  andx  g10457(.a(n11442), .b(n11441), .O(n11443));
  orx   g10458(.a(n11443), .b(n11426), .O(n11444));
  andx  g10459(.a(n11443), .b(n11426), .O(n11445));
  invx  g10460(.a(n11445), .O(n11446));
  andx  g10461(.a(n11446), .b(n11444), .O(n11447));
  orx   g10462(.a(n11447), .b(n11421), .O(n11448));
  andx  g10463(.a(n11447), .b(n11421), .O(n11449));
  invx  g10464(.a(n11449), .O(n11450));
  andx  g10465(.a(n11450), .b(n11448), .O(n11451));
  andx  g10466(.a(n11128), .b(n11081), .O(n11452));
  orx   g10467(.a(n11452), .b(n11125), .O(n11453));
  andx  g10468(.a(n11453), .b(n11451), .O(n11454));
  invx  g10469(.a(n11454), .O(n11455));
  andx  g10470(.a(n11451), .b(n1790), .O(n11456));
  orx   g10471(.a(n11456), .b(n11453), .O(n11457));
  andx  g10472(.a(n11457), .b(n11455), .O(n11458));
  orx   g10473(.a(n11458), .b(n11416), .O(n11459));
  invx  g10474(.a(n11458), .O(n11460));
  orx   g10475(.a(n11460), .b(n11415), .O(n11461));
  andx  g10476(.a(n11461), .b(n11459), .O(po09));
  andx  g10477(.a(n11157), .b(n8062), .O(n11463));
  orx   g10478(.a(n11463), .b(n11161), .O(n11464));
  andx  g10479(.a(n11464), .b(n7982), .O(n11465));
  andx  g10480(.a(n11161), .b(n8062), .O(n11466));
  orx   g10481(.a(n11466), .b(n11465), .O(n11467));
  andx  g10482(.a(n2724), .b(n8062), .O(n11471));
  andx  g10483(.a(n2429), .b(n8131), .O(n11474));
  orx   g10484(.a(n11474), .b(n11471), .O(n11475));
  invx  g10485(.a(n11475), .O(n11477));
  andx  g10486(.a(n8220), .b(n4114), .O(n11480));
  invx  g10487(.a(n11480), .O(n11481));
  orx   g10488(.a(n11173), .b(n11154), .O(n11483));
  andx  g10489(.a(n11483), .b(n11168), .O(n11484));
  orx   g10490(.a(n11484), .b(n11172), .O(n11485));
  andx  g10491(.a(n11485), .b(n11481), .O(n11486));
  invx  g10492(.a(n11172), .O(n11487));
  invx  g10493(.a(n11173), .O(n11488));
  andx  g10494(.a(n11488), .b(n11164), .O(n11489));
  orx   g10495(.a(n11489), .b(n11169), .O(n11490));
  andx  g10496(.a(n11490), .b(n11487), .O(n11491));
  andx  g10497(.a(n11491), .b(n11480), .O(n11492));
  orx   g10498(.a(n11492), .b(n11486), .O(n11493));
  andx  g10499(.a(n11493), .b(n11477), .O(n11494));
  orx   g10500(.a(n11491), .b(n11480), .O(n11496));
  orx   g10501(.a(n11485), .b(n11481), .O(n11497));
  andx  g10502(.a(n11497), .b(n11496), .O(n11498));
  andx  g10503(.a(n11498), .b(n11475), .O(n11499));
  orx   g10504(.a(n11499), .b(n11494), .O(n11500));
  orx   g10505(.a(n11194), .b(n11182), .O(n11501));
  andx  g10506(.a(n11501), .b(n11200), .O(n11502));
  orx   g10507(.a(n11502), .b(n9841), .O(n11503));
  andx  g10508(.a(n11201), .b(n11199), .O(n11504));
  orx   g10509(.a(n11504), .b(n11187), .O(n11505));
  andx  g10510(.a(n8351), .b(n4063), .O(n11506));
  orx   g10511(.a(n11506), .b(n11505), .O(n11507));
  andx  g10512(.a(n11507), .b(n11503), .O(n11508));
  orx   g10513(.a(n11508), .b(n11500), .O(n11509));
  orx   g10514(.a(n11498), .b(n11475), .O(n11510));
  orx   g10515(.a(n11493), .b(n11477), .O(n11511));
  andx  g10516(.a(n11511), .b(n11510), .O(n11512));
  andx  g10517(.a(n11505), .b(n8351), .O(n11513));
  invx  g10518(.a(n11506), .O(n11514));
  andx  g10519(.a(n11514), .b(n11502), .O(n11515));
  orx   g10520(.a(n11515), .b(n11513), .O(n11516));
  orx   g10521(.a(n11516), .b(n11512), .O(n11517));
  andx  g10522(.a(n11517), .b(n11509), .O(n11518));
  andx  g10523(.a(n8603), .b(n3721), .O(n11519));
  andx  g10524(.a(n11211), .b(n11145), .O(n11520));
  invx  g10525(.a(n11520), .O(n11521));
  andx  g10526(.a(n11204), .b(n11140), .O(n11522));
  orx   g10527(.a(n11522), .b(n11142), .O(n11523));
  andx  g10528(.a(n11523), .b(n11521), .O(n11524));
  orx   g10529(.a(n11524), .b(n11519), .O(n11525));
  invx  g10530(.a(n11519), .O(n11526));
  orx   g10531(.a(n11211), .b(n11145), .O(n11527));
  andx  g10532(.a(n11527), .b(n11135), .O(n11528));
  orx   g10533(.a(n11528), .b(n11520), .O(n11529));
  orx   g10534(.a(n11529), .b(n11526), .O(n11530));
  andx  g10535(.a(n11530), .b(n11525), .O(n11531));
  orx   g10536(.a(n11531), .b(n11518), .O(n11532));
  andx  g10537(.a(n11516), .b(n11512), .O(n11533));
  andx  g10538(.a(n11508), .b(n11500), .O(n11534));
  orx   g10539(.a(n11534), .b(n11533), .O(n11535));
  andx  g10540(.a(n11529), .b(n11526), .O(n11536));
  andx  g10541(.a(n11524), .b(n11519), .O(n11537));
  orx   g10542(.a(n11537), .b(n11536), .O(n11538));
  orx   g10543(.a(n11538), .b(n11535), .O(n11539));
  andx  g10544(.a(n11539), .b(n11532), .O(n11540));
  andx  g10545(.a(n11220), .b(n11213), .O(n11541));
  orx   g10546(.a(n11541), .b(n11226), .O(n11542));
  andx  g10547(.a(n11542), .b(n7907), .O(n11543));
  orx   g10548(.a(n11228), .b(n11225), .O(n11544));
  andx  g10549(.a(n11544), .b(n11216), .O(n11545));
  andx  g10550(.a(n7907), .b(n3645), .O(n11546));
  invx  g10551(.a(n11546), .O(n11547));
  andx  g10552(.a(n11547), .b(n11545), .O(n11548));
  orx   g10553(.a(n11548), .b(n11543), .O(n11549));
  andx  g10554(.a(n11549), .b(n11540), .O(n11550));
  andx  g10555(.a(n11538), .b(n11535), .O(n11551));
  andx  g10556(.a(n11531), .b(n11518), .O(n11552));
  orx   g10557(.a(n11552), .b(n11551), .O(n11553));
  orx   g10558(.a(n11545), .b(n10161), .O(n11554));
  orx   g10559(.a(n11546), .b(n11542), .O(n11555));
  andx  g10560(.a(n11555), .b(n11554), .O(n11556));
  andx  g10561(.a(n11556), .b(n11553), .O(n11557));
  orx   g10562(.a(n11557), .b(n11550), .O(n11558));
  andx  g10563(.a(n8852), .b(n3413), .O(n11559));
  invx  g10564(.a(n11559), .O(n11560));
  andx  g10565(.a(n11236), .b(n11231), .O(n11561));
  invx  g10566(.a(n11561), .O(n11562));
  andx  g10567(.a(n11242), .b(n11248), .O(n11563));
  orx   g10568(.a(n11563), .b(n11238), .O(n11564));
  andx  g10569(.a(n11564), .b(n11562), .O(n11565));
  orx   g10570(.a(n11565), .b(n11560), .O(n11566));
  orx   g10571(.a(n11236), .b(n11231), .O(n11567));
  andx  g10572(.a(n11567), .b(n11232), .O(n11568));
  orx   g10573(.a(n11568), .b(n11561), .O(n11569));
  orx   g10574(.a(n11569), .b(n11559), .O(n11570));
  andx  g10575(.a(n11570), .b(n11566), .O(n11571));
  andx  g10576(.a(n11571), .b(n11558), .O(n11572));
  orx   g10577(.a(n11556), .b(n11553), .O(n11573));
  orx   g10578(.a(n11549), .b(n11540), .O(n11574));
  andx  g10579(.a(n11574), .b(n11573), .O(n11575));
  andx  g10580(.a(n11569), .b(n11559), .O(n11576));
  andx  g10581(.a(n11565), .b(n11560), .O(n11577));
  orx   g10582(.a(n11577), .b(n11576), .O(n11578));
  andx  g10583(.a(n11578), .b(n11575), .O(n11579));
  orx   g10584(.a(n11579), .b(n11572), .O(n11580));
  orx   g10585(.a(n11262), .b(n11253), .O(n11581));
  andx  g10586(.a(n11581), .b(n11268), .O(n11582));
  orx   g10587(.a(n11582), .b(n10585), .O(n11583));
  andx  g10588(.a(n11270), .b(n11267), .O(n11584));
  orx   g10589(.a(n11584), .b(n11256), .O(n11585));
  andx  g10590(.a(n9050), .b(n3171), .O(n11586));
  orx   g10591(.a(n11586), .b(n11585), .O(n11587));
  andx  g10592(.a(n11587), .b(n11583), .O(n11588));
  orx   g10593(.a(n11588), .b(n11580), .O(n11589));
  orx   g10594(.a(n11578), .b(n11575), .O(n11590));
  orx   g10595(.a(n11571), .b(n11558), .O(n11591));
  andx  g10596(.a(n11591), .b(n11590), .O(n11592));
  andx  g10597(.a(n11585), .b(n9050), .O(n11593));
  orx   g10598(.a(n10585), .b(n3418), .O(n11594));
  andx  g10599(.a(n11594), .b(n11582), .O(n11595));
  orx   g10600(.a(n11595), .b(n11593), .O(n11596));
  orx   g10601(.a(n11596), .b(n11592), .O(n11597));
  andx  g10602(.a(n11597), .b(n11589), .O(n11598));
  orx   g10603(.a(n9266), .b(n3297), .O(n11599));
  invx  g10604(.a(n11599), .O(n11600));
  orx   g10605(.a(n11284), .b(n11273), .O(n11601));
  andx  g10606(.a(n11284), .b(n11273), .O(n11602));
  orx   g10607(.a(n11602), .b(n11274), .O(n11603));
  andx  g10608(.a(n11603), .b(n11601), .O(n11604));
  orx   g10609(.a(n11604), .b(n11600), .O(n11605));
  andx  g10610(.a(n11278), .b(n11290), .O(n11606));
  orx   g10611(.a(n11278), .b(n11290), .O(n11607));
  andx  g10612(.a(n11607), .b(n11280), .O(n11608));
  orx   g10613(.a(n11608), .b(n11606), .O(n11609));
  orx   g10614(.a(n11609), .b(n11599), .O(n11610));
  andx  g10615(.a(n11610), .b(n11605), .O(n11611));
  orx   g10616(.a(n11611), .b(n11598), .O(n11612));
  andx  g10617(.a(n11596), .b(n11592), .O(n11613));
  andx  g10618(.a(n11588), .b(n11580), .O(n11614));
  orx   g10619(.a(n11614), .b(n11613), .O(n11615));
  andx  g10620(.a(n11609), .b(n11599), .O(n11616));
  andx  g10621(.a(n11604), .b(n11600), .O(n11617));
  orx   g10622(.a(n11617), .b(n11616), .O(n11618));
  orx   g10623(.a(n11618), .b(n11615), .O(n11619));
  andx  g10624(.a(n11619), .b(n11612), .O(n11620));
  andx  g10625(.a(n11303), .b(n11295), .O(n11621));
  orx   g10626(.a(n11621), .b(n11309), .O(n11622));
  andx  g10627(.a(n11622), .b(n9470), .O(n11623));
  orx   g10628(.a(n11310), .b(n11308), .O(n11624));
  andx  g10629(.a(n11624), .b(n11298), .O(n11625));
  andx  g10630(.a(n9470), .b(n3180), .O(n11626));
  invx  g10631(.a(n11626), .O(n11627));
  andx  g10632(.a(n11627), .b(n11625), .O(n11628));
  orx   g10633(.a(n11628), .b(n11623), .O(n11629));
  andx  g10634(.a(n11629), .b(n11620), .O(n11630));
  andx  g10635(.a(n11618), .b(n11615), .O(n11631));
  andx  g10636(.a(n11611), .b(n11598), .O(n11632));
  orx   g10637(.a(n11632), .b(n11631), .O(n11633));
  orx   g10638(.a(n11625), .b(n11012), .O(n11634));
  orx   g10639(.a(n11626), .b(n11622), .O(n11635));
  andx  g10640(.a(n11635), .b(n11634), .O(n11636));
  andx  g10641(.a(n11636), .b(n11633), .O(n11637));
  orx   g10642(.a(n11637), .b(n11630), .O(n11638));
  andx  g10643(.a(n11318), .b(n11313), .O(n11639));
  orx   g10644(.a(n11318), .b(n11313), .O(n11640));
  andx  g10645(.a(n11640), .b(n11314), .O(n11641));
  orx   g10646(.a(n11641), .b(n11639), .O(n11642));
  andx  g10647(.a(n7902), .b(n3284), .O(n11643));
  orx   g10648(.a(n11643), .b(n11642), .O(n11644));
  orx   g10649(.a(n11324), .b(n11330), .O(n11645));
  andx  g10650(.a(n11324), .b(n11330), .O(n11646));
  orx   g10651(.a(n11646), .b(n11320), .O(n11647));
  andx  g10652(.a(n11647), .b(n11645), .O(n11648));
  invx  g10653(.a(n11643), .O(n11649));
  orx   g10654(.a(n11649), .b(n11648), .O(n11650));
  andx  g10655(.a(n11650), .b(n11644), .O(n11651));
  andx  g10656(.a(n11651), .b(n11638), .O(n11652));
  orx   g10657(.a(n11636), .b(n11633), .O(n11653));
  orx   g10658(.a(n11629), .b(n11620), .O(n11654));
  andx  g10659(.a(n11654), .b(n11653), .O(n11655));
  andx  g10660(.a(n11649), .b(n11648), .O(n11656));
  andx  g10661(.a(n11643), .b(n11642), .O(n11657));
  orx   g10662(.a(n11657), .b(n11656), .O(n11658));
  andx  g10663(.a(n11658), .b(n11655), .O(n11659));
  orx   g10664(.a(n11659), .b(n11652), .O(n11660));
  orx   g10665(.a(n11343), .b(n11335), .O(n11661));
  andx  g10666(.a(n11661), .b(n11350), .O(n11662));
  orx   g10667(.a(n11662), .b(n11053), .O(n11663));
  andx  g10668(.a(n11351), .b(n11348), .O(n11664));
  orx   g10669(.a(n11664), .b(n11338), .O(n11665));
  andx  g10670(.a(n10356), .b(n3210), .O(n11666));
  orx   g10671(.a(n11666), .b(n11665), .O(n11667));
  andx  g10672(.a(n11667), .b(n11663), .O(n11668));
  orx   g10673(.a(n11668), .b(n11660), .O(n11669));
  orx   g10674(.a(n11658), .b(n11655), .O(n11670));
  orx   g10675(.a(n11651), .b(n11638), .O(n11671));
  andx  g10676(.a(n11671), .b(n11670), .O(n11672));
  andx  g10677(.a(n11665), .b(n10356), .O(n11673));
  invx  g10678(.a(n11666), .O(n11674));
  andx  g10679(.a(n11674), .b(n11662), .O(n11675));
  orx   g10680(.a(n11675), .b(n11673), .O(n11676));
  orx   g10681(.a(n11676), .b(n11672), .O(n11677));
  andx  g10682(.a(n11677), .b(n11669), .O(n11678));
  orx   g10683(.a(n11367), .b(n11354), .O(n11679));
  andx  g10684(.a(n11367), .b(n11354), .O(n11680));
  orx   g10685(.a(n11680), .b(n11368), .O(n11681));
  andx  g10686(.a(n11681), .b(n11679), .O(n11682));
  andx  g10687(.a(n10751), .b(n3221), .O(n11683));
  invx  g10688(.a(n11683), .O(n11684));
  andx  g10689(.a(n11684), .b(n11682), .O(n11685));
  andx  g10690(.a(n11358), .b(n11374), .O(n11686));
  orx   g10691(.a(n11358), .b(n11374), .O(n11687));
  andx  g10692(.a(n11687), .b(n11359), .O(n11688));
  orx   g10693(.a(n11688), .b(n11686), .O(n11689));
  andx  g10694(.a(n11683), .b(n11689), .O(n11690));
  orx   g10695(.a(n11690), .b(n11685), .O(n11691));
  orx   g10696(.a(n11691), .b(n11678), .O(n11692));
  andx  g10697(.a(n11676), .b(n11672), .O(n11693));
  andx  g10698(.a(n11668), .b(n11660), .O(n11694));
  orx   g10699(.a(n11694), .b(n11693), .O(n11695));
  orx   g10700(.a(n11683), .b(n11689), .O(n11696));
  orx   g10701(.a(n11684), .b(n11682), .O(n11697));
  andx  g10702(.a(n11697), .b(n11696), .O(n11698));
  orx   g10703(.a(n11698), .b(n11695), .O(n11699));
  andx  g10704(.a(n11699), .b(n11692), .O(n11700));
  andx  g10705(.a(n11387), .b(n11379), .O(n11701));
  orx   g10706(.a(n11701), .b(n11393), .O(n11702));
  andx  g10707(.a(n11702), .b(n11120), .O(n11703));
  orx   g10708(.a(n11395), .b(n11392), .O(n11704));
  andx  g10709(.a(n11704), .b(n11383), .O(n11705));
  andx  g10710(.a(n11120), .b(n3230), .O(n11706));
  invx  g10711(.a(n11706), .O(n11707));
  andx  g10712(.a(n11707), .b(n11705), .O(n11708));
  orx   g10713(.a(n11708), .b(n11703), .O(n11709));
  andx  g10714(.a(n11709), .b(n11700), .O(n11710));
  andx  g10715(.a(n11698), .b(n11695), .O(n11711));
  andx  g10716(.a(n11691), .b(n11678), .O(n11712));
  orx   g10717(.a(n11712), .b(n11711), .O(n11713));
  invx  g10718(.a(n11120), .O(n11714));
  orx   g10719(.a(n11705), .b(n11714), .O(n11715));
  orx   g10720(.a(n11706), .b(n11702), .O(n11716));
  andx  g10721(.a(n11716), .b(n11715), .O(n11717));
  andx  g10722(.a(n11717), .b(n11713), .O(n11718));
  orx   g10723(.a(n11718), .b(n11710), .O(n11719));
  andx  g10724(.a(n11409), .b(n11398), .O(n11720));
  invx  g10725(.a(n11720), .O(n11721));
  andx  g10726(.a(n11396), .b(n11392), .O(n11722));
  andx  g10727(.a(n11388), .b(n11379), .O(n11723));
  orx   g10728(.a(n11723), .b(n11722), .O(n11724));
  andx  g10729(.a(n11403), .b(n11724), .O(n11725));
  orx   g10730(.a(n11725), .b(n11405), .O(n11726));
  andx  g10731(.a(n11726), .b(n11721), .O(n11727));
  andx  g10732(.a(n11451), .b(n3258), .O(n11728));
  invx  g10733(.a(n11728), .O(n11729));
  andx  g10734(.a(n11729), .b(n11727), .O(n11730));
  orx   g10735(.a(n11409), .b(n11398), .O(n11731));
  andx  g10736(.a(n11731), .b(n11404), .O(n11732));
  orx   g10737(.a(n11732), .b(n11720), .O(n11733));
  andx  g10738(.a(n11728), .b(n11733), .O(n11734));
  orx   g10739(.a(n11734), .b(n11730), .O(n11735));
  invx  g10740(.a(n11735), .O(n11736));
  andx  g10741(.a(n11736), .b(n11719), .O(n11737));
  orx   g10742(.a(n11717), .b(n11713), .O(n11738));
  orx   g10743(.a(n11709), .b(n11700), .O(n11739));
  andx  g10744(.a(n11739), .b(n11738), .O(n11740));
  andx  g10745(.a(n11735), .b(n11740), .O(n11741));
  orx   g10746(.a(n11741), .b(n11737), .O(n11742));
  invx  g10747(.a(n11121), .O(n11743));
  andx  g10748(.a(n10762), .b(n10693), .O(n11744));
  orx   g10749(.a(n11744), .b(n10758), .O(n11745));
  andx  g10750(.a(n11745), .b(n11743), .O(n11746));
  invx  g10751(.a(n11127), .O(n11747));
  andx  g10752(.a(n11747), .b(n11746), .O(n11748));
  orx   g10753(.a(n11748), .b(n11131), .O(n11749));
  andx  g10754(.a(n11749), .b(n11126), .O(n11750));
  invx  g10755(.a(n11456), .O(n11751));
  andx  g10756(.a(n11751), .b(n11750), .O(n11752));
  orx   g10757(.a(n11752), .b(n11415), .O(n11753));
  andx  g10758(.a(n11753), .b(n11455), .O(n11754));
  andx  g10759(.a(n11754), .b(n11742), .O(n11755));
  invx  g10760(.a(n11742), .O(n11756));
  andx  g10761(.a(n11457), .b(n11416), .O(n11757));
  orx   g10762(.a(n11757), .b(n11454), .O(n11758));
  andx  g10763(.a(n11758), .b(n11756), .O(n11759));
  orx   g10764(.a(n11759), .b(n11755), .O(po10));
  andx  g10765(.a(n8852), .b(n3645), .O(n11761));
  invx  g10766(.a(n11761), .O(n11762));
  orx   g10767(.a(n11548), .b(n11540), .O(n11763));
  andx  g10768(.a(n11763), .b(n11554), .O(n11764));
  andx  g10769(.a(n11764), .b(n11762), .O(n11765));
  andx  g10770(.a(n11555), .b(n11553), .O(n11766));
  orx   g10771(.a(n11766), .b(n11543), .O(n11767));
  andx  g10772(.a(n11767), .b(n8852), .O(n11768));
  orx   g10773(.a(n11768), .b(n11765), .O(n11769));
  andx  g10774(.a(n2429), .b(n8220), .O(n11772));
  andx  g10775(.a(n2724), .b(n8131), .O(n11775));
  orx   g10776(.a(n11775), .b(n11772), .O(n11776));
  andx  g10777(.a(n11157), .b(n8131), .O(n11777));
  orx   g10778(.a(n11777), .b(n11467), .O(n11778));
  andx  g10779(.a(n11778), .b(n8062), .O(n11779));
  andx  g10780(.a(n11467), .b(n8131), .O(n11780));
  orx   g10781(.a(n11780), .b(n11779), .O(n11781));
  invx  g10782(.a(n11781), .O(n11782));
  andx  g10783(.a(n11491), .b(n11477), .O(n11789));
  orx   g10784(.a(n11789), .b(n11481), .O(n11790));
  andx  g10785(.a(n11790), .b(n11490), .O(n11791));
  andx  g10786(.a(n8351), .b(n4114), .O(n11792));
  invx  g10787(.a(n11792), .O(n11793));
  andx  g10788(.a(n11793), .b(n11791), .O(n11794));
  orx   g10789(.a(n11485), .b(n11475), .O(n11795));
  andx  g10790(.a(n11795), .b(n11480), .O(n11796));
  orx   g10791(.a(n11796), .b(n11484), .O(n11797));
  andx  g10792(.a(n11792), .b(n11797), .O(n11798));
  orx   g10793(.a(n11798), .b(n11794), .O(n11799));
  orx   g10794(.a(n11799), .b(n11776), .O(n11800));
  invx  g10795(.a(n11776), .O(n11801));
  orx   g10796(.a(n11792), .b(n11797), .O(n11803));
  orx   g10797(.a(n11793), .b(n11791), .O(n11804));
  andx  g10798(.a(n11804), .b(n11803), .O(n11805));
  orx   g10799(.a(n11805), .b(n11801), .O(n11806));
  andx  g10800(.a(n11806), .b(n11800), .O(n11807));
  andx  g10801(.a(n11507), .b(n11500), .O(n11808));
  orx   g10802(.a(n11808), .b(n11513), .O(n11809));
  andx  g10803(.a(n11809), .b(n8603), .O(n11810));
  orx   g10804(.a(n11515), .b(n11512), .O(n11811));
  andx  g10805(.a(n11811), .b(n11503), .O(n11812));
  andx  g10806(.a(n8603), .b(n4063), .O(n11813));
  invx  g10807(.a(n11813), .O(n11814));
  andx  g10808(.a(n11814), .b(n11812), .O(n11815));
  orx   g10809(.a(n11815), .b(n11810), .O(n11816));
  andx  g10810(.a(n11816), .b(n11807), .O(n11817));
  andx  g10811(.a(n11805), .b(n11801), .O(n11818));
  andx  g10812(.a(n11799), .b(n11776), .O(n11819));
  orx   g10813(.a(n11819), .b(n11818), .O(n11820));
  orx   g10814(.a(n11812), .b(n9680), .O(n11821));
  orx   g10815(.a(n11813), .b(n11809), .O(n11822));
  andx  g10816(.a(n11822), .b(n11821), .O(n11823));
  andx  g10817(.a(n11823), .b(n11820), .O(n11824));
  orx   g10818(.a(n11824), .b(n11817), .O(n11825));
  andx  g10819(.a(n11529), .b(n11518), .O(n11826));
  orx   g10820(.a(n11529), .b(n11518), .O(n11827));
  andx  g10821(.a(n11827), .b(n11519), .O(n11828));
  orx   g10822(.a(n11828), .b(n11826), .O(n11829));
  andx  g10823(.a(n7907), .b(n3721), .O(n11830));
  orx   g10824(.a(n11830), .b(n11829), .O(n11831));
  invx  g10825(.a(n11826), .O(n11832));
  andx  g10826(.a(n11524), .b(n11535), .O(n11833));
  orx   g10827(.a(n11833), .b(n11526), .O(n11834));
  andx  g10828(.a(n11834), .b(n11832), .O(n11835));
  invx  g10829(.a(n11830), .O(n11836));
  orx   g10830(.a(n11836), .b(n11835), .O(n11837));
  andx  g10831(.a(n11837), .b(n11831), .O(n11838));
  andx  g10832(.a(n11838), .b(n11825), .O(n11839));
  orx   g10833(.a(n11823), .b(n11820), .O(n11840));
  orx   g10834(.a(n11816), .b(n11807), .O(n11841));
  andx  g10835(.a(n11841), .b(n11840), .O(n11842));
  andx  g10836(.a(n11836), .b(n11835), .O(n11843));
  andx  g10837(.a(n11830), .b(n11829), .O(n11844));
  orx   g10838(.a(n11844), .b(n11843), .O(n11845));
  andx  g10839(.a(n11845), .b(n11842), .O(n11846));
  orx   g10840(.a(n11846), .b(n11839), .O(n11847));
  andx  g10841(.a(n11847), .b(n11769), .O(n11848));
  orx   g10842(.a(n11767), .b(n11761), .O(n11849));
  orx   g10843(.a(n11764), .b(n11260), .O(n11850));
  andx  g10844(.a(n11850), .b(n11849), .O(n11851));
  orx   g10845(.a(n11845), .b(n11842), .O(n11852));
  orx   g10846(.a(n11838), .b(n11825), .O(n11853));
  andx  g10847(.a(n11853), .b(n11852), .O(n11854));
  andx  g10848(.a(n11854), .b(n11851), .O(n11855));
  orx   g10849(.a(n11855), .b(n11848), .O(n11856));
  andx  g10850(.a(n9050), .b(n3413), .O(n11857));
  andx  g10851(.a(n11569), .b(n11575), .O(n11858));
  orx   g10852(.a(n11569), .b(n11575), .O(n11859));
  andx  g10853(.a(n11859), .b(n11559), .O(n11860));
  orx   g10854(.a(n11860), .b(n11858), .O(n11861));
  andx  g10855(.a(n11861), .b(n11857), .O(n11862));
  invx  g10856(.a(n11857), .O(n11863));
  invx  g10857(.a(n11858), .O(n11864));
  andx  g10858(.a(n11565), .b(n11558), .O(n11865));
  orx   g10859(.a(n11865), .b(n11560), .O(n11866));
  andx  g10860(.a(n11866), .b(n11864), .O(n11867));
  andx  g10861(.a(n11867), .b(n11863), .O(n11868));
  orx   g10862(.a(n11868), .b(n11862), .O(n11869));
  orx   g10863(.a(n11869), .b(n11856), .O(n11870));
  orx   g10864(.a(n11854), .b(n11851), .O(n11871));
  orx   g10865(.a(n11847), .b(n11769), .O(n11872));
  andx  g10866(.a(n11872), .b(n11871), .O(n11873));
  orx   g10867(.a(n11867), .b(n11863), .O(n11874));
  orx   g10868(.a(n11861), .b(n11857), .O(n11875));
  andx  g10869(.a(n11875), .b(n11874), .O(n11876));
  orx   g10870(.a(n11876), .b(n11873), .O(n11877));
  andx  g10871(.a(n11877), .b(n11870), .O(n11878));
  andx  g10872(.a(n11587), .b(n11580), .O(n11879));
  orx   g10873(.a(n11879), .b(n11593), .O(n11880));
  andx  g10874(.a(n11880), .b(n9267), .O(n11881));
  orx   g10875(.a(n11595), .b(n11592), .O(n11882));
  andx  g10876(.a(n11882), .b(n11583), .O(n11883));
  andx  g10877(.a(n9267), .b(n3171), .O(n11884));
  invx  g10878(.a(n11884), .O(n11885));
  andx  g10879(.a(n11885), .b(n11883), .O(n11886));
  orx   g10880(.a(n11886), .b(n11881), .O(n11887));
  andx  g10881(.a(n11887), .b(n11878), .O(n11888));
  andx  g10882(.a(n11876), .b(n11873), .O(n11889));
  andx  g10883(.a(n11869), .b(n11856), .O(n11890));
  orx   g10884(.a(n11890), .b(n11889), .O(n11891));
  orx   g10885(.a(n11883), .b(n9266), .O(n11892));
  orx   g10886(.a(n11884), .b(n11880), .O(n11893));
  andx  g10887(.a(n11893), .b(n11892), .O(n11894));
  andx  g10888(.a(n11894), .b(n11891), .O(n11895));
  orx   g10889(.a(n11895), .b(n11888), .O(n11896));
  andx  g10890(.a(n9470), .b(n3429), .O(n11897));
  invx  g10891(.a(n11897), .O(n11898));
  andx  g10892(.a(n11609), .b(n11598), .O(n11899));
  orx   g10893(.a(n11609), .b(n11598), .O(n11900));
  andx  g10894(.a(n11900), .b(n11600), .O(n11901));
  orx   g10895(.a(n11901), .b(n11899), .O(n11902));
  andx  g10896(.a(n11902), .b(n11898), .O(n11903));
  invx  g10897(.a(n11899), .O(n11904));
  andx  g10898(.a(n11604), .b(n11615), .O(n11905));
  orx   g10899(.a(n11905), .b(n11599), .O(n11906));
  andx  g10900(.a(n11906), .b(n11904), .O(n11907));
  andx  g10901(.a(n11907), .b(n11897), .O(n11908));
  orx   g10902(.a(n11908), .b(n11903), .O(n11909));
  andx  g10903(.a(n11909), .b(n11896), .O(n11910));
  orx   g10904(.a(n11894), .b(n11891), .O(n11911));
  orx   g10905(.a(n11887), .b(n11878), .O(n11912));
  andx  g10906(.a(n11912), .b(n11911), .O(n11913));
  orx   g10907(.a(n11907), .b(n11897), .O(n11914));
  orx   g10908(.a(n11902), .b(n11898), .O(n11915));
  andx  g10909(.a(n11915), .b(n11914), .O(n11916));
  andx  g10910(.a(n11916), .b(n11913), .O(n11917));
  orx   g10911(.a(n11917), .b(n11910), .O(n11918));
  orx   g10912(.a(n11628), .b(n11620), .O(n11919));
  andx  g10913(.a(n11919), .b(n11634), .O(n11920));
  orx   g10914(.a(n11920), .b(n11349), .O(n11921));
  andx  g10915(.a(n11635), .b(n11633), .O(n11922));
  orx   g10916(.a(n11922), .b(n11623), .O(n11923));
  andx  g10917(.a(n7902), .b(n3180), .O(n11924));
  orx   g10918(.a(n11924), .b(n11923), .O(n11925));
  andx  g10919(.a(n11925), .b(n11921), .O(n11926));
  orx   g10920(.a(n11926), .b(n11918), .O(n11927));
  orx   g10921(.a(n11916), .b(n11913), .O(n11928));
  orx   g10922(.a(n11909), .b(n11896), .O(n11929));
  andx  g10923(.a(n11929), .b(n11928), .O(n11930));
  andx  g10924(.a(n11923), .b(n7902), .O(n11931));
  invx  g10925(.a(n11924), .O(n11932));
  andx  g10926(.a(n11932), .b(n11920), .O(n11933));
  orx   g10927(.a(n11933), .b(n11931), .O(n11934));
  orx   g10928(.a(n11934), .b(n11930), .O(n11935));
  andx  g10929(.a(n11935), .b(n11927), .O(n11936));
  orx   g10930(.a(n11648), .b(n11638), .O(n11937));
  andx  g10931(.a(n11648), .b(n11638), .O(n11938));
  orx   g10932(.a(n11938), .b(n11649), .O(n11939));
  andx  g10933(.a(n11939), .b(n11937), .O(n11940));
  andx  g10934(.a(n10356), .b(n3284), .O(n11941));
  invx  g10935(.a(n11941), .O(n11942));
  andx  g10936(.a(n11942), .b(n11940), .O(n11943));
  andx  g10937(.a(n11642), .b(n11655), .O(n11944));
  orx   g10938(.a(n11642), .b(n11655), .O(n11945));
  andx  g10939(.a(n11945), .b(n11643), .O(n11946));
  orx   g10940(.a(n11946), .b(n11944), .O(n11947));
  andx  g10941(.a(n11941), .b(n11947), .O(n11948));
  orx   g10942(.a(n11948), .b(n11943), .O(n11949));
  orx   g10943(.a(n11949), .b(n11936), .O(n11950));
  andx  g10944(.a(n11934), .b(n11930), .O(n11951));
  andx  g10945(.a(n11926), .b(n11918), .O(n11952));
  orx   g10946(.a(n11952), .b(n11951), .O(n11953));
  orx   g10947(.a(n11941), .b(n11947), .O(n11954));
  orx   g10948(.a(n11942), .b(n11940), .O(n11955));
  andx  g10949(.a(n11955), .b(n11954), .O(n11956));
  orx   g10950(.a(n11956), .b(n11953), .O(n11957));
  andx  g10951(.a(n11957), .b(n11950), .O(n11958));
  andx  g10952(.a(n11667), .b(n11660), .O(n11959));
  orx   g10953(.a(n11959), .b(n11673), .O(n11960));
  andx  g10954(.a(n11960), .b(n10751), .O(n11961));
  orx   g10955(.a(n11675), .b(n11672), .O(n11962));
  andx  g10956(.a(n11962), .b(n11663), .O(n11963));
  andx  g10957(.a(n10751), .b(n3210), .O(n11964));
  invx  g10958(.a(n11964), .O(n11965));
  andx  g10959(.a(n11965), .b(n11963), .O(n11966));
  orx   g10960(.a(n11966), .b(n11961), .O(n11967));
  andx  g10961(.a(n11967), .b(n11958), .O(n11968));
  andx  g10962(.a(n11956), .b(n11953), .O(n11969));
  andx  g10963(.a(n11949), .b(n11936), .O(n11970));
  orx   g10964(.a(n11970), .b(n11969), .O(n11971));
  orx   g10965(.a(n11963), .b(n11380), .O(n11972));
  orx   g10966(.a(n11964), .b(n11960), .O(n11973));
  andx  g10967(.a(n11973), .b(n11972), .O(n11974));
  andx  g10968(.a(n11974), .b(n11971), .O(n11975));
  orx   g10969(.a(n11975), .b(n11968), .O(n11976));
  andx  g10970(.a(n11689), .b(n11678), .O(n11977));
  orx   g10971(.a(n11689), .b(n11678), .O(n11978));
  andx  g10972(.a(n11978), .b(n11683), .O(n11979));
  orx   g10973(.a(n11979), .b(n11977), .O(n11980));
  andx  g10974(.a(n11120), .b(n3221), .O(n11981));
  orx   g10975(.a(n11981), .b(n11980), .O(n11982));
  orx   g10976(.a(n11682), .b(n11695), .O(n11983));
  andx  g10977(.a(n11682), .b(n11695), .O(n11984));
  orx   g10978(.a(n11984), .b(n11684), .O(n11985));
  andx  g10979(.a(n11985), .b(n11983), .O(n11986));
  invx  g10980(.a(n11981), .O(n11987));
  orx   g10981(.a(n11987), .b(n11986), .O(n11988));
  andx  g10982(.a(n11988), .b(n11982), .O(n11989));
  andx  g10983(.a(n11989), .b(n11976), .O(n11990));
  orx   g10984(.a(n11974), .b(n11971), .O(n11991));
  orx   g10985(.a(n11967), .b(n11958), .O(n11992));
  andx  g10986(.a(n11992), .b(n11991), .O(n11993));
  andx  g10987(.a(n11987), .b(n11986), .O(n11994));
  andx  g10988(.a(n11981), .b(n11980), .O(n11995));
  orx   g10989(.a(n11995), .b(n11994), .O(n11996));
  andx  g10990(.a(n11996), .b(n11993), .O(n11997));
  orx   g10991(.a(n11997), .b(n11990), .O(n11998));
  invx  g10992(.a(n11448), .O(n11999));
  orx   g10993(.a(n11449), .b(n11999), .O(n12000));
  orx   g10994(.a(n11708), .b(n11700), .O(n12001));
  andx  g10995(.a(n12001), .b(n11715), .O(n12002));
  orx   g10996(.a(n12002), .b(n12000), .O(n12003));
  andx  g10997(.a(n11716), .b(n11713), .O(n12004));
  orx   g10998(.a(n12004), .b(n11703), .O(n12005));
  andx  g10999(.a(n11451), .b(n3230), .O(n12006));
  orx   g11000(.a(n12006), .b(n12005), .O(n12007));
  andx  g11001(.a(n12007), .b(n12003), .O(n12008));
  orx   g11002(.a(n12008), .b(n11998), .O(n12009));
  orx   g11003(.a(n11996), .b(n11993), .O(n12010));
  orx   g11004(.a(n11989), .b(n11976), .O(n12011));
  andx  g11005(.a(n12011), .b(n12010), .O(n12012));
  andx  g11006(.a(n12005), .b(n11451), .O(n12013));
  invx  g11007(.a(n12006), .O(n12014));
  andx  g11008(.a(n12014), .b(n12002), .O(n12015));
  orx   g11009(.a(n12015), .b(n12013), .O(n12016));
  orx   g11010(.a(n12016), .b(n12012), .O(n12017));
  andx  g11011(.a(n12017), .b(n12009), .O(n12018));
  andx  g11012(.a(n11728), .b(n11740), .O(n12019));
  andx  g11013(.a(n11733), .b(n11740), .O(n12020));
  orx   g11014(.a(n12020), .b(n11734), .O(n12021));
  orx   g11015(.a(n12021), .b(n12019), .O(n12022));
  andx  g11016(.a(n12022), .b(n12018), .O(n12023));
  orx   g11017(.a(n12023), .b(n11754), .O(n12024));
  andx  g11018(.a(n12016), .b(n12012), .O(n12025));
  andx  g11019(.a(n12008), .b(n11998), .O(n12026));
  orx   g11020(.a(n12026), .b(n12025), .O(n12027));
  invx  g11021(.a(n12019), .O(n12028));
  orx   g11022(.a(n11729), .b(n11727), .O(n12029));
  orx   g11023(.a(n11727), .b(n11719), .O(n12030));
  andx  g11024(.a(n12030), .b(n12029), .O(n12031));
  andx  g11025(.a(n12031), .b(n12028), .O(n12032));
  andx  g11026(.a(n12032), .b(n12027), .O(n12033));
  orx   g11027(.a(n12033), .b(n11756), .O(n12034));
  orx   g11028(.a(n12034), .b(n12024), .O(n12035));
  andx  g11029(.a(n11758), .b(n11742), .O(n12036));
  andx  g11030(.a(n12022), .b(n12027), .O(n12037));
  andx  g11031(.a(n12032), .b(n12018), .O(n12038));
  orx   g11032(.a(n12038), .b(n12037), .O(n12039));
  orx   g11033(.a(n12039), .b(n12036), .O(n12040));
  andx  g11034(.a(n12040), .b(n12035), .O(po11));
  orx   g11035(.a(n12032), .b(n12027), .O(n12042));
  orx   g11036(.a(n12015), .b(n12012), .O(n12043));
  andx  g11037(.a(n12043), .b(n12003), .O(n12044));
  andx  g11038(.a(n9050), .b(n3645), .O(n12045));
  invx  g11039(.a(n12045), .O(n12046));
  orx   g11040(.a(n11854), .b(n11765), .O(n12047));
  andx  g11041(.a(n12047), .b(n11850), .O(n12048));
  andx  g11042(.a(n12048), .b(n12046), .O(n12049));
  andx  g11043(.a(n11847), .b(n11849), .O(n12050));
  orx   g11044(.a(n12050), .b(n11768), .O(n12051));
  andx  g11045(.a(n12051), .b(n9050), .O(n12052));
  orx   g11046(.a(n12052), .b(n12049), .O(n12053));
  andx  g11047(.a(n2724), .b(n8220), .O(n12056));
  andx  g11048(.a(n2429), .b(n8351), .O(n12059));
  orx   g11049(.a(n12059), .b(n12056), .O(n12060));
  andx  g11050(.a(n11157), .b(n8220), .O(n12061));
  invx  g11051(.a(n12061), .O(n12062));
  andx  g11052(.a(n12062), .b(n11782), .O(n12063));
  orx   g11053(.a(n12063), .b(n8770), .O(n12064));
  andx  g11054(.a(n11781), .b(n8220), .O(n12065));
  invx  g11055(.a(n12065), .O(n12066));
  andx  g11056(.a(n12066), .b(n12064), .O(n12067));
  invx  g11057(.a(n12060), .O(n12069));
  andx  g11058(.a(n11791), .b(n11801), .O(n12075));
  orx   g11059(.a(n12075), .b(n11793), .O(n12076));
  andx  g11060(.a(n12076), .b(n11790), .O(n12077));
  andx  g11061(.a(n8603), .b(n4114), .O(n12078));
  invx  g11062(.a(n12078), .O(n12079));
  andx  g11063(.a(n12079), .b(n12077), .O(n12080));
  orx   g11064(.a(n11797), .b(n11776), .O(n12081));
  andx  g11065(.a(n12081), .b(n11792), .O(n12082));
  orx   g11066(.a(n12082), .b(n11796), .O(n12083));
  andx  g11067(.a(n12078), .b(n12083), .O(n12084));
  orx   g11068(.a(n12084), .b(n12080), .O(n12085));
  orx   g11069(.a(n12085), .b(n12060), .O(n12086));
  orx   g11070(.a(n12078), .b(n12083), .O(n12087));
  orx   g11071(.a(n12079), .b(n12077), .O(n12088));
  andx  g11072(.a(n12088), .b(n12087), .O(n12089));
  orx   g11073(.a(n12089), .b(n12069), .O(n12090));
  andx  g11074(.a(n12090), .b(n12086), .O(n12091));
  andx  g11075(.a(n11822), .b(n11820), .O(n12092));
  orx   g11076(.a(n12092), .b(n11810), .O(n12093));
  andx  g11077(.a(n12093), .b(n7907), .O(n12094));
  orx   g11078(.a(n11815), .b(n11807), .O(n12095));
  andx  g11079(.a(n12095), .b(n11821), .O(n12096));
  andx  g11080(.a(n7907), .b(n4063), .O(n12097));
  invx  g11081(.a(n12097), .O(n12098));
  andx  g11082(.a(n12098), .b(n12096), .O(n12099));
  orx   g11083(.a(n12099), .b(n12094), .O(n12100));
  andx  g11084(.a(n12100), .b(n12091), .O(n12101));
  andx  g11085(.a(n12089), .b(n12069), .O(n12102));
  andx  g11086(.a(n12085), .b(n12060), .O(n12103));
  orx   g11087(.a(n12103), .b(n12102), .O(n12104));
  orx   g11088(.a(n12096), .b(n10161), .O(n12105));
  orx   g11089(.a(n12097), .b(n12093), .O(n12106));
  andx  g11090(.a(n12106), .b(n12105), .O(n12107));
  andx  g11091(.a(n12107), .b(n12104), .O(n12108));
  orx   g11092(.a(n12108), .b(n12101), .O(n12109));
  andx  g11093(.a(n11829), .b(n11842), .O(n12110));
  orx   g11094(.a(n11829), .b(n11842), .O(n12111));
  andx  g11095(.a(n12111), .b(n11830), .O(n12112));
  orx   g11096(.a(n12112), .b(n12110), .O(n12113));
  andx  g11097(.a(n8852), .b(n3721), .O(n12114));
  orx   g11098(.a(n12114), .b(n12113), .O(n12115));
  invx  g11099(.a(n12110), .O(n12116));
  andx  g11100(.a(n11835), .b(n11825), .O(n12117));
  orx   g11101(.a(n12117), .b(n11836), .O(n12118));
  andx  g11102(.a(n12118), .b(n12116), .O(n12119));
  invx  g11103(.a(n12114), .O(n12120));
  orx   g11104(.a(n12120), .b(n12119), .O(n12121));
  andx  g11105(.a(n12121), .b(n12115), .O(n12122));
  andx  g11106(.a(n12122), .b(n12109), .O(n12123));
  orx   g11107(.a(n12107), .b(n12104), .O(n12124));
  orx   g11108(.a(n12100), .b(n12091), .O(n12125));
  andx  g11109(.a(n12125), .b(n12124), .O(n12126));
  andx  g11110(.a(n12120), .b(n12119), .O(n12127));
  andx  g11111(.a(n12114), .b(n12113), .O(n12128));
  orx   g11112(.a(n12128), .b(n12127), .O(n12129));
  andx  g11113(.a(n12129), .b(n12126), .O(n12130));
  orx   g11114(.a(n12130), .b(n12123), .O(n12131));
  andx  g11115(.a(n12131), .b(n12053), .O(n12132));
  orx   g11116(.a(n12051), .b(n12045), .O(n12133));
  orx   g11117(.a(n12048), .b(n10585), .O(n12134));
  andx  g11118(.a(n12134), .b(n12133), .O(n12135));
  orx   g11119(.a(n12129), .b(n12126), .O(n12136));
  orx   g11120(.a(n12122), .b(n12109), .O(n12137));
  andx  g11121(.a(n12137), .b(n12136), .O(n12138));
  andx  g11122(.a(n12138), .b(n12135), .O(n12139));
  orx   g11123(.a(n12139), .b(n12132), .O(n12140));
  andx  g11124(.a(n9267), .b(n3413), .O(n12141));
  andx  g11125(.a(n11861), .b(n11856), .O(n12142));
  invx  g11126(.a(n12142), .O(n12143));
  andx  g11127(.a(n11867), .b(n11873), .O(n12144));
  orx   g11128(.a(n12144), .b(n11863), .O(n12145));
  andx  g11129(.a(n12145), .b(n12143), .O(n12146));
  orx   g11130(.a(n12146), .b(n12141), .O(n12147));
  invx  g11131(.a(n12141), .O(n12148));
  orx   g11132(.a(n11861), .b(n11856), .O(n12149));
  andx  g11133(.a(n12149), .b(n11857), .O(n12150));
  orx   g11134(.a(n12150), .b(n12142), .O(n12151));
  orx   g11135(.a(n12151), .b(n12148), .O(n12152));
  andx  g11136(.a(n12152), .b(n12147), .O(n12153));
  orx   g11137(.a(n12153), .b(n12140), .O(n12154));
  orx   g11138(.a(n12138), .b(n12135), .O(n12155));
  orx   g11139(.a(n12131), .b(n12053), .O(n12156));
  andx  g11140(.a(n12156), .b(n12155), .O(n12157));
  andx  g11141(.a(n12151), .b(n12148), .O(n12158));
  andx  g11142(.a(n12146), .b(n12141), .O(n12159));
  orx   g11143(.a(n12159), .b(n12158), .O(n12160));
  orx   g11144(.a(n12160), .b(n12157), .O(n12161));
  andx  g11145(.a(n12161), .b(n12154), .O(n12162));
  andx  g11146(.a(n11893), .b(n11891), .O(n12163));
  orx   g11147(.a(n12163), .b(n11881), .O(n12164));
  andx  g11148(.a(n12164), .b(n9470), .O(n12165));
  andx  g11149(.a(n9470), .b(n3171), .O(n12166));
  orx   g11150(.a(n12166), .b(n12164), .O(n12167));
  invx  g11151(.a(n12167), .O(n12168));
  orx   g11152(.a(n12168), .b(n12165), .O(n12169));
  andx  g11153(.a(n12169), .b(n12162), .O(n12170));
  andx  g11154(.a(n12160), .b(n12157), .O(n12171));
  andx  g11155(.a(n12153), .b(n12140), .O(n12172));
  orx   g11156(.a(n12172), .b(n12171), .O(n12173));
  invx  g11157(.a(n12165), .O(n12174));
  andx  g11158(.a(n12167), .b(n12174), .O(n12175));
  andx  g11159(.a(n12175), .b(n12173), .O(n12176));
  orx   g11160(.a(n12176), .b(n12170), .O(n12177));
  andx  g11161(.a(n7902), .b(n3429), .O(n12178));
  invx  g11162(.a(n12178), .O(n12179));
  andx  g11163(.a(n11902), .b(n11913), .O(n12180));
  orx   g11164(.a(n11902), .b(n11913), .O(n12181));
  andx  g11165(.a(n12181), .b(n11897), .O(n12182));
  orx   g11166(.a(n12182), .b(n12180), .O(n12183));
  andx  g11167(.a(n12183), .b(n12179), .O(n12184));
  invx  g11168(.a(n12180), .O(n12185));
  andx  g11169(.a(n11907), .b(n11896), .O(n12186));
  orx   g11170(.a(n12186), .b(n11898), .O(n12187));
  andx  g11171(.a(n12187), .b(n12185), .O(n12188));
  andx  g11172(.a(n12188), .b(n12178), .O(n12189));
  orx   g11173(.a(n12189), .b(n12184), .O(n12190));
  andx  g11174(.a(n12190), .b(n12177), .O(n12191));
  orx   g11175(.a(n12175), .b(n12173), .O(n12192));
  orx   g11176(.a(n12169), .b(n12162), .O(n12193));
  andx  g11177(.a(n12193), .b(n12192), .O(n12194));
  orx   g11178(.a(n12188), .b(n12178), .O(n12195));
  orx   g11179(.a(n12183), .b(n12179), .O(n12196));
  andx  g11180(.a(n12196), .b(n12195), .O(n12197));
  andx  g11181(.a(n12197), .b(n12194), .O(n12198));
  orx   g11182(.a(n12198), .b(n12191), .O(n12199));
  orx   g11183(.a(n11933), .b(n11930), .O(n12200));
  andx  g11184(.a(n12200), .b(n11921), .O(n12201));
  orx   g11185(.a(n12201), .b(n11053), .O(n12202));
  andx  g11186(.a(n11925), .b(n11918), .O(n12203));
  orx   g11187(.a(n12203), .b(n11931), .O(n12204));
  andx  g11188(.a(n10356), .b(n3180), .O(n12205));
  orx   g11189(.a(n12205), .b(n12204), .O(n12206));
  andx  g11190(.a(n12206), .b(n12202), .O(n12207));
  orx   g11191(.a(n12207), .b(n12199), .O(n12208));
  orx   g11192(.a(n12197), .b(n12194), .O(n12209));
  orx   g11193(.a(n12190), .b(n12177), .O(n12210));
  andx  g11194(.a(n12210), .b(n12209), .O(n12211));
  andx  g11195(.a(n12204), .b(n10356), .O(n12212));
  invx  g11196(.a(n12205), .O(n12213));
  andx  g11197(.a(n12213), .b(n12201), .O(n12214));
  orx   g11198(.a(n12214), .b(n12212), .O(n12215));
  orx   g11199(.a(n12215), .b(n12211), .O(n12216));
  andx  g11200(.a(n12216), .b(n12208), .O(n12217));
  orx   g11201(.a(n11940), .b(n11953), .O(n12218));
  andx  g11202(.a(n11940), .b(n11953), .O(n12219));
  orx   g11203(.a(n12219), .b(n11942), .O(n12220));
  andx  g11204(.a(n12220), .b(n12218), .O(n12221));
  andx  g11205(.a(n10751), .b(n3284), .O(n12222));
  invx  g11206(.a(n12222), .O(n12223));
  andx  g11207(.a(n12223), .b(n12221), .O(n12224));
  andx  g11208(.a(n11947), .b(n11936), .O(n12225));
  orx   g11209(.a(n11947), .b(n11936), .O(n12226));
  andx  g11210(.a(n12226), .b(n11941), .O(n12227));
  orx   g11211(.a(n12227), .b(n12225), .O(n12228));
  andx  g11212(.a(n12222), .b(n12228), .O(n12229));
  orx   g11213(.a(n12229), .b(n12224), .O(n12230));
  orx   g11214(.a(n12230), .b(n12217), .O(n12231));
  andx  g11215(.a(n12215), .b(n12211), .O(n12232));
  andx  g11216(.a(n12207), .b(n12199), .O(n12233));
  orx   g11217(.a(n12233), .b(n12232), .O(n12234));
  orx   g11218(.a(n12222), .b(n12228), .O(n12235));
  orx   g11219(.a(n12223), .b(n12221), .O(n12236));
  andx  g11220(.a(n12236), .b(n12235), .O(n12237));
  orx   g11221(.a(n12237), .b(n12234), .O(n12238));
  andx  g11222(.a(n12238), .b(n12231), .O(n12239));
  andx  g11223(.a(n11973), .b(n11971), .O(n12240));
  orx   g11224(.a(n12240), .b(n11961), .O(n12241));
  andx  g11225(.a(n12241), .b(n11120), .O(n12242));
  orx   g11226(.a(n11966), .b(n11958), .O(n12243));
  andx  g11227(.a(n12243), .b(n11972), .O(n12244));
  andx  g11228(.a(n11120), .b(n3210), .O(n12245));
  invx  g11229(.a(n12245), .O(n12246));
  andx  g11230(.a(n12246), .b(n12244), .O(n12247));
  orx   g11231(.a(n12247), .b(n12242), .O(n12248));
  andx  g11232(.a(n12248), .b(n12239), .O(n12249));
  andx  g11233(.a(n12237), .b(n12234), .O(n12250));
  andx  g11234(.a(n12230), .b(n12217), .O(n12251));
  orx   g11235(.a(n12251), .b(n12250), .O(n12252));
  orx   g11236(.a(n12244), .b(n11714), .O(n12253));
  orx   g11237(.a(n12245), .b(n12241), .O(n12254));
  andx  g11238(.a(n12254), .b(n12253), .O(n12255));
  andx  g11239(.a(n12255), .b(n12252), .O(n12256));
  orx   g11240(.a(n12256), .b(n12249), .O(n12257));
  orx   g11241(.a(n11986), .b(n11976), .O(n12258));
  andx  g11242(.a(n11986), .b(n11976), .O(n12259));
  orx   g11243(.a(n12259), .b(n11987), .O(n12260));
  andx  g11244(.a(n12260), .b(n12258), .O(n12261));
  andx  g11245(.a(n11451), .b(n3221), .O(n12262));
  invx  g11246(.a(n12262), .O(n12263));
  andx  g11247(.a(n12263), .b(n12261), .O(n12264));
  andx  g11248(.a(n11980), .b(n11993), .O(n12265));
  orx   g11249(.a(n11980), .b(n11993), .O(n12266));
  andx  g11250(.a(n12266), .b(n11981), .O(n12267));
  orx   g11251(.a(n12267), .b(n12265), .O(n12268));
  andx  g11252(.a(n12262), .b(n12268), .O(n12269));
  orx   g11253(.a(n12269), .b(n12264), .O(n12270));
  orx   g11254(.a(n12270), .b(n12257), .O(n12271));
  orx   g11255(.a(n12255), .b(n12252), .O(n12272));
  orx   g11256(.a(n12248), .b(n12239), .O(n12273));
  andx  g11257(.a(n12273), .b(n12272), .O(n12274));
  orx   g11258(.a(n12262), .b(n12268), .O(n12275));
  orx   g11259(.a(n12263), .b(n12261), .O(n12276));
  andx  g11260(.a(n12276), .b(n12275), .O(n12277));
  orx   g11261(.a(n12277), .b(n12274), .O(n12278));
  andx  g11262(.a(n12278), .b(n12271), .O(n12279));
  andx  g11263(.a(n12279), .b(n12044), .O(n12280));
  andx  g11264(.a(n12007), .b(n11998), .O(n12281));
  orx   g11265(.a(n12281), .b(n12013), .O(n12282));
  andx  g11266(.a(n12277), .b(n12274), .O(n12283));
  andx  g11267(.a(n12270), .b(n12257), .O(n12284));
  orx   g11268(.a(n12284), .b(n12283), .O(n12285));
  andx  g11269(.a(n12285), .b(n12282), .O(n12286));
  orx   g11270(.a(n12286), .b(n12280), .O(n12287));
  andx  g11271(.a(n12287), .b(n12042), .O(n12288));
  andx  g11272(.a(n12288), .b(n12035), .O(n12289));
  orx   g11273(.a(n12285), .b(n12282), .O(n12290));
  orx   g11274(.a(n12279), .b(n12044), .O(n12291));
  andx  g11275(.a(n12291), .b(n12290), .O(n12292));
  andx  g11276(.a(n12292), .b(n12023), .O(n12293));
  andx  g11277(.a(n12042), .b(n11758), .O(n12294));
  invx  g11278(.a(n12034), .O(n12295));
  andx  g11279(.a(n12295), .b(n12294), .O(n12296));
  andx  g11280(.a(n12292), .b(n12296), .O(n12297));
  orx   g11281(.a(n12297), .b(n12293), .O(n12298));
  orx   g11282(.a(n12298), .b(n12289), .O(po12));
  andx  g11283(.a(n12035), .b(n12042), .O(n12300));
  orx   g11284(.a(n12300), .b(n12292), .O(n12301));
  invx  g11285(.a(n12301), .O(n12302));
  andx  g11286(.a(n12262), .b(n12274), .O(n12303));
  orx   g11287(.a(n12262), .b(n12274), .O(n12304));
  andx  g11288(.a(n12304), .b(n12268), .O(n12305));
  orx   g11289(.a(n12305), .b(n12303), .O(n12306));
  andx  g11290(.a(n12254), .b(n12252), .O(n12307));
  orx   g11291(.a(n12307), .b(n12242), .O(n12308));
  andx  g11292(.a(n11451), .b(n3210), .O(n12309));
  orx   g11293(.a(n12309), .b(n12308), .O(n12310));
  orx   g11294(.a(n12247), .b(n12239), .O(n12311));
  andx  g11295(.a(n12311), .b(n12253), .O(n12312));
  orx   g11296(.a(n12312), .b(n12000), .O(n12313));
  andx  g11297(.a(n12313), .b(n12310), .O(n12314));
  andx  g11298(.a(n9267), .b(n3645), .O(n12315));
  invx  g11299(.a(n12315), .O(n12316));
  orx   g11300(.a(n12138), .b(n12049), .O(n12317));
  andx  g11301(.a(n12317), .b(n12134), .O(n12318));
  andx  g11302(.a(n12318), .b(n12316), .O(n12319));
  andx  g11303(.a(n12131), .b(n12133), .O(n12320));
  orx   g11304(.a(n12320), .b(n12052), .O(n12321));
  andx  g11305(.a(n12321), .b(n9267), .O(n12322));
  orx   g11306(.a(n12322), .b(n12319), .O(n12323));
  andx  g11307(.a(n8852), .b(n4063), .O(n12324));
  andx  g11308(.a(n12106), .b(n12104), .O(n12325));
  orx   g11309(.a(n12325), .b(n12094), .O(n12326));
  orx   g11310(.a(n12326), .b(n12324), .O(n12327));
  orx   g11311(.a(n12099), .b(n12091), .O(n12328));
  andx  g11312(.a(n12328), .b(n12105), .O(n12329));
  orx   g11313(.a(n12329), .b(n11260), .O(n12330));
  andx  g11314(.a(n12330), .b(n12327), .O(n12331));
  andx  g11315(.a(n12067), .b(n12062), .O(n12332));
  orx   g11316(.a(n12332), .b(n9841), .O(n12333));
  orx   g11317(.a(n12067), .b(n8675), .O(n12334));
  andx  g11318(.a(n12334), .b(n12333), .O(n12335));
  andx  g11319(.a(n2724), .b(n8351), .O(n12338));
  andx  g11320(.a(n2429), .b(n8603), .O(n12341));
  orx   g11321(.a(n12341), .b(n12338), .O(n12342));
  invx  g11322(.a(n12342), .O(n12344));
  andx  g11323(.a(n7907), .b(n4114), .O(n12348));
  andx  g11324(.a(n12077), .b(n12069), .O(n12350));
  orx   g11325(.a(n12350), .b(n12079), .O(n12351));
  invx  g11326(.a(n12351), .O(n12352));
  orx   g11327(.a(n12352), .b(n12082), .O(n12353));
  andx  g11328(.a(n12353), .b(n12348), .O(n12354));
  invx  g11329(.a(n12348), .O(n12355));
  andx  g11330(.a(n12351), .b(n12076), .O(n12357));
  andx  g11331(.a(n12357), .b(n12355), .O(n12358));
  orx   g11332(.a(n12358), .b(n12354), .O(n12359));
  orx   g11333(.a(n12359), .b(n12342), .O(n12360));
  orx   g11334(.a(n12357), .b(n12355), .O(n12361));
  orx   g11335(.a(n12353), .b(n12348), .O(n12362));
  andx  g11336(.a(n12362), .b(n12361), .O(n12363));
  orx   g11337(.a(n12363), .b(n12344), .O(n12364));
  andx  g11338(.a(n12364), .b(n12360), .O(n12365));
  orx   g11339(.a(n12365), .b(n12331), .O(n12366));
  invx  g11340(.a(n12324), .O(n12367));
  andx  g11341(.a(n12329), .b(n12367), .O(n12368));
  andx  g11342(.a(n12326), .b(n8852), .O(n12369));
  orx   g11343(.a(n12369), .b(n12368), .O(n12370));
  andx  g11344(.a(n12363), .b(n12344), .O(n12371));
  andx  g11345(.a(n12359), .b(n12342), .O(n12372));
  orx   g11346(.a(n12372), .b(n12371), .O(n12373));
  orx   g11347(.a(n12373), .b(n12370), .O(n12374));
  andx  g11348(.a(n12374), .b(n12366), .O(n12375));
  andx  g11349(.a(n12113), .b(n12126), .O(n12376));
  orx   g11350(.a(n12113), .b(n12126), .O(n12377));
  andx  g11351(.a(n12377), .b(n12114), .O(n12378));
  orx   g11352(.a(n12378), .b(n12376), .O(n12379));
  andx  g11353(.a(n9050), .b(n3721), .O(n12380));
  orx   g11354(.a(n12380), .b(n12379), .O(n12381));
  invx  g11355(.a(n12376), .O(n12382));
  andx  g11356(.a(n12119), .b(n12109), .O(n12383));
  orx   g11357(.a(n12383), .b(n12120), .O(n12384));
  andx  g11358(.a(n12384), .b(n12382), .O(n12385));
  invx  g11359(.a(n12380), .O(n12386));
  orx   g11360(.a(n12386), .b(n12385), .O(n12387));
  andx  g11361(.a(n12387), .b(n12381), .O(n12388));
  andx  g11362(.a(n12388), .b(n12375), .O(n12389));
  andx  g11363(.a(n12373), .b(n12370), .O(n12390));
  andx  g11364(.a(n12365), .b(n12331), .O(n12391));
  orx   g11365(.a(n12391), .b(n12390), .O(n12392));
  andx  g11366(.a(n12386), .b(n12385), .O(n12393));
  andx  g11367(.a(n12380), .b(n12379), .O(n12394));
  orx   g11368(.a(n12394), .b(n12393), .O(n12395));
  andx  g11369(.a(n12395), .b(n12392), .O(n12396));
  orx   g11370(.a(n12396), .b(n12389), .O(n12397));
  andx  g11371(.a(n12397), .b(n12323), .O(n12398));
  orx   g11372(.a(n12321), .b(n12315), .O(n12399));
  orx   g11373(.a(n12318), .b(n9266), .O(n12400));
  andx  g11374(.a(n12400), .b(n12399), .O(n12401));
  orx   g11375(.a(n12395), .b(n12392), .O(n12402));
  orx   g11376(.a(n12388), .b(n12375), .O(n12403));
  andx  g11377(.a(n12403), .b(n12402), .O(n12404));
  andx  g11378(.a(n12404), .b(n12401), .O(n12405));
  orx   g11379(.a(n12405), .b(n12398), .O(n12406));
  andx  g11380(.a(n9470), .b(n3413), .O(n12407));
  andx  g11381(.a(n12151), .b(n12140), .O(n12408));
  invx  g11382(.a(n12408), .O(n12409));
  andx  g11383(.a(n12146), .b(n12157), .O(n12410));
  orx   g11384(.a(n12410), .b(n12148), .O(n12411));
  andx  g11385(.a(n12411), .b(n12409), .O(n12412));
  orx   g11386(.a(n12412), .b(n12407), .O(n12413));
  invx  g11387(.a(n12407), .O(n12414));
  orx   g11388(.a(n12151), .b(n12140), .O(n12415));
  andx  g11389(.a(n12415), .b(n12141), .O(n12416));
  orx   g11390(.a(n12416), .b(n12408), .O(n12417));
  orx   g11391(.a(n12417), .b(n12414), .O(n12418));
  andx  g11392(.a(n12418), .b(n12413), .O(n12419));
  orx   g11393(.a(n12419), .b(n12406), .O(n12420));
  orx   g11394(.a(n12404), .b(n12401), .O(n12421));
  orx   g11395(.a(n12397), .b(n12323), .O(n12422));
  andx  g11396(.a(n12422), .b(n12421), .O(n12423));
  andx  g11397(.a(n12417), .b(n12414), .O(n12424));
  andx  g11398(.a(n12412), .b(n12407), .O(n12425));
  orx   g11399(.a(n12425), .b(n12424), .O(n12426));
  orx   g11400(.a(n12426), .b(n12423), .O(n12427));
  andx  g11401(.a(n12427), .b(n12420), .O(n12428));
  andx  g11402(.a(n12167), .b(n12173), .O(n12429));
  orx   g11403(.a(n12429), .b(n12165), .O(n12430));
  andx  g11404(.a(n12430), .b(n7902), .O(n12431));
  orx   g11405(.a(n12168), .b(n12162), .O(n12432));
  andx  g11406(.a(n12432), .b(n12174), .O(n12433));
  andx  g11407(.a(n7902), .b(n3171), .O(n12434));
  invx  g11408(.a(n12434), .O(n12435));
  andx  g11409(.a(n12435), .b(n12433), .O(n12436));
  orx   g11410(.a(n12436), .b(n12431), .O(n12437));
  andx  g11411(.a(n12437), .b(n12428), .O(n12438));
  andx  g11412(.a(n12426), .b(n12423), .O(n12439));
  andx  g11413(.a(n12419), .b(n12406), .O(n12440));
  orx   g11414(.a(n12440), .b(n12439), .O(n12441));
  orx   g11415(.a(n12433), .b(n11349), .O(n12442));
  orx   g11416(.a(n12434), .b(n12430), .O(n12443));
  andx  g11417(.a(n12443), .b(n12442), .O(n12444));
  andx  g11418(.a(n12444), .b(n12441), .O(n12445));
  orx   g11419(.a(n12445), .b(n12438), .O(n12446));
  andx  g11420(.a(n10356), .b(n3429), .O(n12447));
  invx  g11421(.a(n12447), .O(n12448));
  andx  g11422(.a(n12183), .b(n12194), .O(n12449));
  orx   g11423(.a(n12183), .b(n12194), .O(n12450));
  andx  g11424(.a(n12450), .b(n12178), .O(n12451));
  orx   g11425(.a(n12451), .b(n12449), .O(n12452));
  andx  g11426(.a(n12452), .b(n12448), .O(n12453));
  invx  g11427(.a(n12449), .O(n12454));
  andx  g11428(.a(n12188), .b(n12177), .O(n12455));
  orx   g11429(.a(n12455), .b(n12179), .O(n12456));
  andx  g11430(.a(n12456), .b(n12454), .O(n12457));
  andx  g11431(.a(n12457), .b(n12447), .O(n12458));
  orx   g11432(.a(n12458), .b(n12453), .O(n12459));
  andx  g11433(.a(n12459), .b(n12446), .O(n12460));
  orx   g11434(.a(n12444), .b(n12441), .O(n12461));
  orx   g11435(.a(n12437), .b(n12428), .O(n12462));
  andx  g11436(.a(n12462), .b(n12461), .O(n12463));
  orx   g11437(.a(n12457), .b(n12447), .O(n12464));
  orx   g11438(.a(n12452), .b(n12448), .O(n12465));
  andx  g11439(.a(n12465), .b(n12464), .O(n12466));
  andx  g11440(.a(n12466), .b(n12463), .O(n12467));
  orx   g11441(.a(n12467), .b(n12460), .O(n12468));
  andx  g11442(.a(n12206), .b(n12199), .O(n12469));
  orx   g11443(.a(n12469), .b(n12212), .O(n12470));
  andx  g11444(.a(n12470), .b(n10751), .O(n12471));
  invx  g11445(.a(n12471), .O(n12472));
  andx  g11446(.a(n10751), .b(n3180), .O(n12473));
  orx   g11447(.a(n12473), .b(n12470), .O(n12474));
  andx  g11448(.a(n12474), .b(n12472), .O(n12475));
  orx   g11449(.a(n12475), .b(n12468), .O(n12476));
  orx   g11450(.a(n12466), .b(n12463), .O(n12477));
  orx   g11451(.a(n12459), .b(n12446), .O(n12478));
  andx  g11452(.a(n12478), .b(n12477), .O(n12479));
  invx  g11453(.a(n12474), .O(n12480));
  orx   g11454(.a(n12480), .b(n12471), .O(n12481));
  orx   g11455(.a(n12481), .b(n12479), .O(n12482));
  andx  g11456(.a(n12482), .b(n12476), .O(n12483));
  andx  g11457(.a(n12228), .b(n12217), .O(n12484));
  invx  g11458(.a(n12484), .O(n12485));
  andx  g11459(.a(n12221), .b(n12234), .O(n12486));
  orx   g11460(.a(n12486), .b(n12223), .O(n12487));
  andx  g11461(.a(n12487), .b(n12485), .O(n12488));
  andx  g11462(.a(n11120), .b(n3284), .O(n12489));
  invx  g11463(.a(n12489), .O(n12490));
  andx  g11464(.a(n12490), .b(n12488), .O(n12491));
  orx   g11465(.a(n12228), .b(n12217), .O(n12492));
  andx  g11466(.a(n12492), .b(n12222), .O(n12493));
  orx   g11467(.a(n12493), .b(n12484), .O(n12494));
  andx  g11468(.a(n12489), .b(n12494), .O(n12495));
  orx   g11469(.a(n12495), .b(n12491), .O(n12496));
  orx   g11470(.a(n12496), .b(n12483), .O(n12497));
  andx  g11471(.a(n12481), .b(n12479), .O(n12498));
  andx  g11472(.a(n12475), .b(n12468), .O(n12499));
  orx   g11473(.a(n12499), .b(n12498), .O(n12500));
  orx   g11474(.a(n12489), .b(n12494), .O(n12501));
  orx   g11475(.a(n12490), .b(n12488), .O(n12502));
  andx  g11476(.a(n12502), .b(n12501), .O(n12503));
  orx   g11477(.a(n12503), .b(n12500), .O(n12504));
  andx  g11478(.a(n12504), .b(n12497), .O(n12505));
  orx   g11479(.a(n12505), .b(n12314), .O(n12506));
  orx   g11480(.a(n12000), .b(n3270), .O(n12507));
  andx  g11481(.a(n12507), .b(n12312), .O(n12508));
  andx  g11482(.a(n12308), .b(n11451), .O(n12509));
  orx   g11483(.a(n12509), .b(n12508), .O(n12510));
  andx  g11484(.a(n12503), .b(n12500), .O(n12511));
  andx  g11485(.a(n12496), .b(n12483), .O(n12512));
  orx   g11486(.a(n12512), .b(n12511), .O(n12513));
  orx   g11487(.a(n12513), .b(n12510), .O(n12514));
  andx  g11488(.a(n12514), .b(n12506), .O(n12515));
  andx  g11489(.a(n12515), .b(n12306), .O(n12516));
  orx   g11490(.a(n12263), .b(n12257), .O(n12517));
  andx  g11491(.a(n12263), .b(n12257), .O(n12518));
  orx   g11492(.a(n12518), .b(n12261), .O(n12519));
  andx  g11493(.a(n12519), .b(n12517), .O(n12520));
  andx  g11494(.a(n12513), .b(n12510), .O(n12521));
  andx  g11495(.a(n12505), .b(n12314), .O(n12522));
  orx   g11496(.a(n12522), .b(n12521), .O(n12523));
  andx  g11497(.a(n12523), .b(n12520), .O(n12524));
  orx   g11498(.a(n12524), .b(n12516), .O(n12525));
  andx  g11499(.a(n12279), .b(n12282), .O(n12526));
  orx   g11500(.a(n12526), .b(n12525), .O(n12527));
  andx  g11501(.a(n12526), .b(n12525), .O(n12528));
  invx  g11502(.a(n12528), .O(n12529));
  andx  g11503(.a(n12529), .b(n12527), .O(n12530));
  orx   g11504(.a(n12530), .b(n12302), .O(n12531));
  invx  g11505(.a(n12530), .O(n12532));
  orx   g11506(.a(n12532), .b(n12301), .O(n12533));
  andx  g11507(.a(n12533), .b(n12531), .O(po13));
  andx  g11508(.a(n12523), .b(n12306), .O(n12535));
  invx  g11509(.a(n12535), .O(n12536));
  andx  g11510(.a(n12513), .b(n12310), .O(n12537));
  orx   g11511(.a(n12537), .b(n12509), .O(n12538));
  invx  g11512(.a(n12538), .O(n12539));
  andx  g11513(.a(n9470), .b(n3645), .O(n12540));
  invx  g11514(.a(n12540), .O(n12541));
  orx   g11515(.a(n12404), .b(n12319), .O(n12542));
  andx  g11516(.a(n12542), .b(n12400), .O(n12543));
  andx  g11517(.a(n12543), .b(n12541), .O(n12544));
  andx  g11518(.a(n12397), .b(n12399), .O(n12545));
  orx   g11519(.a(n12545), .b(n12322), .O(n12546));
  andx  g11520(.a(n12546), .b(n9470), .O(n12547));
  orx   g11521(.a(n12547), .b(n12544), .O(n12548));
  andx  g11522(.a(n9050), .b(n4063), .O(n12549));
  andx  g11523(.a(n12373), .b(n12327), .O(n12550));
  orx   g11524(.a(n12550), .b(n12369), .O(n12551));
  orx   g11525(.a(n12551), .b(n12549), .O(n12552));
  orx   g11526(.a(n12365), .b(n12368), .O(n12553));
  andx  g11527(.a(n12553), .b(n12330), .O(n12554));
  orx   g11528(.a(n12554), .b(n10585), .O(n12555));
  andx  g11529(.a(n12555), .b(n12552), .O(n12556));
  andx  g11530(.a(n2429), .b(n7907), .O(n12559));
  andx  g11531(.a(n2724), .b(n8603), .O(n12562));
  orx   g11532(.a(n12562), .b(n12559), .O(n12563));
  invx  g11533(.a(n12335), .O(n12564));
  andx  g11534(.a(n11157), .b(n8603), .O(n12565));
  orx   g11535(.a(n12565), .b(n12564), .O(n12566));
  andx  g11536(.a(n12566), .b(n8351), .O(n12567));
  andx  g11537(.a(n12564), .b(n8603), .O(n12568));
  orx   g11538(.a(n12568), .b(n12567), .O(n12569));
  invx  g11539(.a(n12563), .O(n12572));
  andx  g11540(.a(n12357), .b(n12344), .O(n12578));
  orx   g11541(.a(n12578), .b(n12355), .O(n12579));
  andx  g11542(.a(n12579), .b(n12351), .O(n12580));
  andx  g11543(.a(n8852), .b(n4114), .O(n12581));
  invx  g11544(.a(n12581), .O(n12582));
  andx  g11545(.a(n12582), .b(n12580), .O(n12583));
  invx  g11546(.a(n12579), .O(n12584));
  orx   g11547(.a(n12584), .b(n12352), .O(n12585));
  andx  g11548(.a(n12581), .b(n12585), .O(n12586));
  orx   g11549(.a(n12586), .b(n12583), .O(n12587));
  orx   g11550(.a(n12587), .b(n12563), .O(n12588));
  orx   g11551(.a(n12581), .b(n12585), .O(n12589));
  orx   g11552(.a(n12582), .b(n12580), .O(n12590));
  andx  g11553(.a(n12590), .b(n12589), .O(n12591));
  orx   g11554(.a(n12591), .b(n12572), .O(n12592));
  andx  g11555(.a(n12592), .b(n12588), .O(n12593));
  orx   g11556(.a(n12593), .b(n12556), .O(n12594));
  invx  g11557(.a(n12549), .O(n12595));
  andx  g11558(.a(n12554), .b(n12595), .O(n12596));
  andx  g11559(.a(n12551), .b(n9050), .O(n12597));
  orx   g11560(.a(n12597), .b(n12596), .O(n12598));
  andx  g11561(.a(n12591), .b(n12572), .O(n12599));
  andx  g11562(.a(n12587), .b(n12563), .O(n12600));
  orx   g11563(.a(n12600), .b(n12599), .O(n12601));
  orx   g11564(.a(n12601), .b(n12598), .O(n12602));
  andx  g11565(.a(n12602), .b(n12594), .O(n12603));
  andx  g11566(.a(n12379), .b(n12392), .O(n12604));
  orx   g11567(.a(n12379), .b(n12392), .O(n12605));
  andx  g11568(.a(n12605), .b(n12380), .O(n12606));
  orx   g11569(.a(n12606), .b(n12604), .O(n12607));
  andx  g11570(.a(n9267), .b(n3721), .O(n12608));
  orx   g11571(.a(n12608), .b(n12607), .O(n12609));
  invx  g11572(.a(n12604), .O(n12610));
  andx  g11573(.a(n12385), .b(n12375), .O(n12611));
  orx   g11574(.a(n12611), .b(n12386), .O(n12612));
  andx  g11575(.a(n12612), .b(n12610), .O(n12613));
  invx  g11576(.a(n12608), .O(n12614));
  orx   g11577(.a(n12614), .b(n12613), .O(n12615));
  andx  g11578(.a(n12615), .b(n12609), .O(n12616));
  andx  g11579(.a(n12616), .b(n12603), .O(n12617));
  andx  g11580(.a(n12601), .b(n12598), .O(n12618));
  andx  g11581(.a(n12593), .b(n12556), .O(n12619));
  orx   g11582(.a(n12619), .b(n12618), .O(n12620));
  andx  g11583(.a(n12614), .b(n12613), .O(n12621));
  andx  g11584(.a(n12608), .b(n12607), .O(n12622));
  orx   g11585(.a(n12622), .b(n12621), .O(n12623));
  andx  g11586(.a(n12623), .b(n12620), .O(n12624));
  orx   g11587(.a(n12624), .b(n12617), .O(n12625));
  andx  g11588(.a(n12625), .b(n12548), .O(n12626));
  orx   g11589(.a(n12546), .b(n12540), .O(n12627));
  orx   g11590(.a(n12543), .b(n11012), .O(n12628));
  andx  g11591(.a(n12628), .b(n12627), .O(n12629));
  orx   g11592(.a(n12623), .b(n12620), .O(n12630));
  orx   g11593(.a(n12616), .b(n12603), .O(n12631));
  andx  g11594(.a(n12631), .b(n12630), .O(n12632));
  andx  g11595(.a(n12632), .b(n12629), .O(n12633));
  orx   g11596(.a(n12633), .b(n12626), .O(n12634));
  andx  g11597(.a(n7902), .b(n3413), .O(n12635));
  andx  g11598(.a(n12417), .b(n12406), .O(n12636));
  invx  g11599(.a(n12636), .O(n12637));
  andx  g11600(.a(n12412), .b(n12423), .O(n12638));
  orx   g11601(.a(n12638), .b(n12414), .O(n12639));
  andx  g11602(.a(n12639), .b(n12637), .O(n12640));
  orx   g11603(.a(n12640), .b(n12635), .O(n12641));
  invx  g11604(.a(n12635), .O(n12642));
  orx   g11605(.a(n12417), .b(n12406), .O(n12643));
  andx  g11606(.a(n12643), .b(n12407), .O(n12644));
  orx   g11607(.a(n12644), .b(n12636), .O(n12645));
  orx   g11608(.a(n12645), .b(n12642), .O(n12646));
  andx  g11609(.a(n12646), .b(n12641), .O(n12647));
  orx   g11610(.a(n12647), .b(n12634), .O(n12648));
  orx   g11611(.a(n12632), .b(n12629), .O(n12649));
  orx   g11612(.a(n12625), .b(n12548), .O(n12650));
  andx  g11613(.a(n12650), .b(n12649), .O(n12651));
  andx  g11614(.a(n12645), .b(n12642), .O(n12652));
  andx  g11615(.a(n12640), .b(n12635), .O(n12653));
  orx   g11616(.a(n12653), .b(n12652), .O(n12654));
  orx   g11617(.a(n12654), .b(n12651), .O(n12655));
  andx  g11618(.a(n12655), .b(n12648), .O(n12656));
  andx  g11619(.a(n12443), .b(n12441), .O(n12657));
  orx   g11620(.a(n12657), .b(n12431), .O(n12658));
  andx  g11621(.a(n12658), .b(n10356), .O(n12659));
  orx   g11622(.a(n12436), .b(n12428), .O(n12660));
  andx  g11623(.a(n12660), .b(n12442), .O(n12661));
  andx  g11624(.a(n10356), .b(n3171), .O(n12662));
  invx  g11625(.a(n12662), .O(n12663));
  andx  g11626(.a(n12663), .b(n12661), .O(n12664));
  orx   g11627(.a(n12664), .b(n12659), .O(n12665));
  andx  g11628(.a(n12665), .b(n12656), .O(n12666));
  andx  g11629(.a(n12654), .b(n12651), .O(n12667));
  andx  g11630(.a(n12647), .b(n12634), .O(n12668));
  orx   g11631(.a(n12668), .b(n12667), .O(n12669));
  orx   g11632(.a(n12661), .b(n11053), .O(n12670));
  orx   g11633(.a(n12662), .b(n12658), .O(n12671));
  andx  g11634(.a(n12671), .b(n12670), .O(n12672));
  andx  g11635(.a(n12672), .b(n12669), .O(n12673));
  orx   g11636(.a(n12673), .b(n12666), .O(n12674));
  andx  g11637(.a(n10751), .b(n3429), .O(n12675));
  invx  g11638(.a(n12675), .O(n12676));
  andx  g11639(.a(n12452), .b(n12463), .O(n12677));
  orx   g11640(.a(n12452), .b(n12463), .O(n12678));
  andx  g11641(.a(n12678), .b(n12447), .O(n12679));
  orx   g11642(.a(n12679), .b(n12677), .O(n12680));
  andx  g11643(.a(n12680), .b(n12676), .O(n12681));
  invx  g11644(.a(n12677), .O(n12682));
  andx  g11645(.a(n12457), .b(n12446), .O(n12683));
  orx   g11646(.a(n12683), .b(n12448), .O(n12684));
  andx  g11647(.a(n12684), .b(n12682), .O(n12685));
  andx  g11648(.a(n12685), .b(n12675), .O(n12686));
  orx   g11649(.a(n12686), .b(n12681), .O(n12687));
  andx  g11650(.a(n12687), .b(n12674), .O(n12688));
  invx  g11651(.a(n12688), .O(n12689));
  orx   g11652(.a(n12687), .b(n12674), .O(n12690));
  andx  g11653(.a(n12690), .b(n12689), .O(n12691));
  andx  g11654(.a(n12474), .b(n12468), .O(n12692));
  orx   g11655(.a(n12692), .b(n12471), .O(n12693));
  andx  g11656(.a(n12693), .b(n11120), .O(n12694));
  andx  g11657(.a(n11120), .b(n3180), .O(n12695));
  orx   g11658(.a(n12695), .b(n12693), .O(n12696));
  invx  g11659(.a(n12696), .O(n12697));
  orx   g11660(.a(n12697), .b(n12694), .O(n12698));
  andx  g11661(.a(n12698), .b(n12691), .O(n12699));
  invx  g11662(.a(n12690), .O(n12700));
  orx   g11663(.a(n12700), .b(n12688), .O(n12701));
  invx  g11664(.a(n12694), .O(n12702));
  andx  g11665(.a(n12696), .b(n12702), .O(n12703));
  andx  g11666(.a(n12703), .b(n12701), .O(n12704));
  orx   g11667(.a(n12704), .b(n12699), .O(n12705));
  andx  g11668(.a(n12494), .b(n12483), .O(n12706));
  orx   g11669(.a(n12494), .b(n12483), .O(n12707));
  andx  g11670(.a(n12707), .b(n12489), .O(n12708));
  orx   g11671(.a(n12708), .b(n12706), .O(n12709));
  andx  g11672(.a(n11451), .b(n3284), .O(n12710));
  orx   g11673(.a(n12710), .b(n12709), .O(n12711));
  invx  g11674(.a(n12706), .O(n12712));
  andx  g11675(.a(n12488), .b(n12500), .O(n12713));
  orx   g11676(.a(n12713), .b(n12490), .O(n12714));
  andx  g11677(.a(n12714), .b(n12712), .O(n12715));
  invx  g11678(.a(n12710), .O(n12716));
  orx   g11679(.a(n12716), .b(n12715), .O(n12717));
  andx  g11680(.a(n12717), .b(n12711), .O(n12718));
  andx  g11681(.a(n12718), .b(n12705), .O(n12719));
  orx   g11682(.a(n12703), .b(n12701), .O(n12720));
  orx   g11683(.a(n12698), .b(n12691), .O(n12721));
  andx  g11684(.a(n12721), .b(n12720), .O(n12722));
  andx  g11685(.a(n12716), .b(n12715), .O(n12723));
  andx  g11686(.a(n12710), .b(n12709), .O(n12724));
  orx   g11687(.a(n12724), .b(n12723), .O(n12725));
  andx  g11688(.a(n12725), .b(n12722), .O(n12726));
  orx   g11689(.a(n12726), .b(n12719), .O(n12727));
  orx   g11690(.a(n12727), .b(n12539), .O(n12728));
  orx   g11691(.a(n12725), .b(n12722), .O(n12729));
  orx   g11692(.a(n12718), .b(n12705), .O(n12730));
  andx  g11693(.a(n12730), .b(n12729), .O(n12731));
  orx   g11694(.a(n12731), .b(n12538), .O(n12732));
  andx  g11695(.a(n12732), .b(n12728), .O(n12733));
  orx   g11696(.a(n12733), .b(n12536), .O(n12734));
  andx  g11697(.a(n12731), .b(n12538), .O(n12735));
  andx  g11698(.a(n12727), .b(n12539), .O(n12736));
  orx   g11699(.a(n12736), .b(n12735), .O(n12737));
  orx   g11700(.a(n12737), .b(n12535), .O(n12738));
  andx  g11701(.a(n12738), .b(n12734), .O(n12739));
  invx  g11702(.a(n12739), .O(n12740));
  andx  g11703(.a(n12527), .b(n12302), .O(n12741));
  orx   g11704(.a(n12741), .b(n12528), .O(n12742));
  andx  g11705(.a(n12742), .b(n12740), .O(n12743));
  invx  g11706(.a(n12742), .O(n12744));
  andx  g11707(.a(n12744), .b(n12739), .O(n12745));
  orx   g11708(.a(n12745), .b(n12743), .O(po14));
  andx  g11709(.a(n7902), .b(n3645), .O(n12747));
  invx  g11710(.a(n12747), .O(n12748));
  orx   g11711(.a(n12632), .b(n12544), .O(n12749));
  andx  g11712(.a(n12749), .b(n12628), .O(n12750));
  andx  g11713(.a(n12750), .b(n12748), .O(n12751));
  andx  g11714(.a(n12625), .b(n12627), .O(n12752));
  orx   g11715(.a(n12752), .b(n12547), .O(n12753));
  andx  g11716(.a(n12753), .b(n7902), .O(n12754));
  orx   g11717(.a(n12754), .b(n12751), .O(n12755));
  andx  g11718(.a(n9267), .b(n4063), .O(n12756));
  andx  g11719(.a(n12601), .b(n12552), .O(n12757));
  orx   g11720(.a(n12757), .b(n12597), .O(n12758));
  orx   g11721(.a(n12758), .b(n12756), .O(n12759));
  orx   g11722(.a(n12593), .b(n12596), .O(n12760));
  andx  g11723(.a(n12760), .b(n12555), .O(n12761));
  orx   g11724(.a(n12761), .b(n9266), .O(n12762));
  andx  g11725(.a(n12762), .b(n12759), .O(n12763));
  andx  g11726(.a(n11157), .b(n7907), .O(n12764));
  orx   g11727(.a(n12764), .b(n12569), .O(n12765));
  andx  g11728(.a(n12765), .b(n8603), .O(n12766));
  andx  g11729(.a(n12569), .b(n7907), .O(n12767));
  orx   g11730(.a(n12767), .b(n12766), .O(n12768));
  invx  g11731(.a(n12768), .O(n12769));
  andx  g11732(.a(n9050), .b(n4114), .O(n12782));
  invx  g11733(.a(n12782), .O(n12783));
  andx  g11734(.a(n12580), .b(n12572), .O(n12786));
  orx   g11735(.a(n12786), .b(n12582), .O(n12787));
  andx  g11736(.a(n12787), .b(n12579), .O(n12788));
  orx   g11737(.a(n12788), .b(n12783), .O(n12789));
  invx  g11738(.a(n12789), .O(n12790));
  andx  g11739(.a(n12788), .b(n12783), .O(n12791));
  orx   g11740(.a(n12791), .b(n12790), .O(n12792));
  orx   g11741(.a(n12792), .b(n8852), .O(n12793));
  invx  g11742(.a(n12791), .O(n12794));
  andx  g11743(.a(n12794), .b(n12789), .O(n12795));
  orx   g11744(.a(n12795), .b(n11260), .O(n12796));
  andx  g11745(.a(n12796), .b(n12793), .O(n12797));
  orx   g11746(.a(n12797), .b(n12763), .O(n12798));
  invx  g11747(.a(n12756), .O(n12799));
  andx  g11748(.a(n12761), .b(n12799), .O(n12800));
  andx  g11749(.a(n12758), .b(n9267), .O(n12801));
  orx   g11750(.a(n12801), .b(n12800), .O(n12802));
  andx  g11751(.a(n12795), .b(n11260), .O(n12803));
  andx  g11752(.a(n12792), .b(n8852), .O(n12804));
  orx   g11753(.a(n12804), .b(n12803), .O(n12805));
  orx   g11754(.a(n12805), .b(n12802), .O(n12806));
  andx  g11755(.a(n12806), .b(n12798), .O(n12807));
  andx  g11756(.a(n12607), .b(n12620), .O(n12808));
  orx   g11757(.a(n12607), .b(n12620), .O(n12809));
  andx  g11758(.a(n12809), .b(n12608), .O(n12810));
  orx   g11759(.a(n12810), .b(n12808), .O(n12811));
  andx  g11760(.a(n9470), .b(n3721), .O(n12812));
  orx   g11761(.a(n12812), .b(n12811), .O(n12813));
  invx  g11762(.a(n12808), .O(n12814));
  andx  g11763(.a(n12613), .b(n12603), .O(n12815));
  orx   g11764(.a(n12815), .b(n12614), .O(n12816));
  andx  g11765(.a(n12816), .b(n12814), .O(n12817));
  invx  g11766(.a(n12812), .O(n12818));
  orx   g11767(.a(n12818), .b(n12817), .O(n12819));
  andx  g11768(.a(n12819), .b(n12813), .O(n12820));
  andx  g11769(.a(n12820), .b(n12807), .O(n12821));
  andx  g11770(.a(n12805), .b(n12802), .O(n12822));
  andx  g11771(.a(n12797), .b(n12763), .O(n12823));
  orx   g11772(.a(n12823), .b(n12822), .O(n12824));
  andx  g11773(.a(n12818), .b(n12817), .O(n12825));
  andx  g11774(.a(n12812), .b(n12811), .O(n12826));
  orx   g11775(.a(n12826), .b(n12825), .O(n12827));
  andx  g11776(.a(n12827), .b(n12824), .O(n12828));
  orx   g11777(.a(n12828), .b(n12821), .O(n12829));
  andx  g11778(.a(n12829), .b(n12755), .O(n12830));
  orx   g11779(.a(n12753), .b(n12747), .O(n12831));
  orx   g11780(.a(n12750), .b(n11349), .O(n12832));
  andx  g11781(.a(n12832), .b(n12831), .O(n12833));
  orx   g11782(.a(n12827), .b(n12824), .O(n12834));
  orx   g11783(.a(n12820), .b(n12807), .O(n12835));
  andx  g11784(.a(n12835), .b(n12834), .O(n12836));
  andx  g11785(.a(n12836), .b(n12833), .O(n12837));
  orx   g11786(.a(n12837), .b(n12830), .O(n12838));
  andx  g11787(.a(n10356), .b(n3413), .O(n12839));
  andx  g11788(.a(n12645), .b(n12634), .O(n12840));
  invx  g11789(.a(n12840), .O(n12841));
  andx  g11790(.a(n12640), .b(n12651), .O(n12842));
  orx   g11791(.a(n12842), .b(n12642), .O(n12843));
  andx  g11792(.a(n12843), .b(n12841), .O(n12844));
  orx   g11793(.a(n12844), .b(n12839), .O(n12845));
  invx  g11794(.a(n12839), .O(n12846));
  orx   g11795(.a(n12645), .b(n12634), .O(n12847));
  andx  g11796(.a(n12847), .b(n12635), .O(n12848));
  orx   g11797(.a(n12848), .b(n12840), .O(n12849));
  orx   g11798(.a(n12849), .b(n12846), .O(n12850));
  andx  g11799(.a(n12850), .b(n12845), .O(n12851));
  orx   g11800(.a(n12851), .b(n12838), .O(n12852));
  orx   g11801(.a(n12836), .b(n12833), .O(n12853));
  orx   g11802(.a(n12829), .b(n12755), .O(n12854));
  andx  g11803(.a(n12854), .b(n12853), .O(n12855));
  andx  g11804(.a(n12849), .b(n12846), .O(n12856));
  andx  g11805(.a(n12844), .b(n12839), .O(n12857));
  orx   g11806(.a(n12857), .b(n12856), .O(n12858));
  orx   g11807(.a(n12858), .b(n12855), .O(n12859));
  andx  g11808(.a(n12859), .b(n12852), .O(n12860));
  andx  g11809(.a(n12671), .b(n12669), .O(n12861));
  orx   g11810(.a(n12861), .b(n12659), .O(n12862));
  andx  g11811(.a(n12862), .b(n10751), .O(n12863));
  orx   g11812(.a(n12664), .b(n12656), .O(n12864));
  andx  g11813(.a(n12864), .b(n12670), .O(n12865));
  andx  g11814(.a(n10751), .b(n3171), .O(n12866));
  invx  g11815(.a(n12866), .O(n12867));
  andx  g11816(.a(n12867), .b(n12865), .O(n12868));
  orx   g11817(.a(n12868), .b(n12863), .O(n12869));
  andx  g11818(.a(n12869), .b(n12860), .O(n12870));
  andx  g11819(.a(n12858), .b(n12855), .O(n12871));
  andx  g11820(.a(n12851), .b(n12838), .O(n12872));
  orx   g11821(.a(n12872), .b(n12871), .O(n12873));
  orx   g11822(.a(n12865), .b(n11380), .O(n12874));
  orx   g11823(.a(n12866), .b(n12862), .O(n12875));
  andx  g11824(.a(n12875), .b(n12874), .O(n12876));
  andx  g11825(.a(n12876), .b(n12873), .O(n12877));
  orx   g11826(.a(n12877), .b(n12870), .O(n12878));
  andx  g11827(.a(n11120), .b(n3429), .O(n12879));
  invx  g11828(.a(n12879), .O(n12880));
  orx   g11829(.a(n12672), .b(n12669), .O(n12881));
  orx   g11830(.a(n12665), .b(n12656), .O(n12882));
  andx  g11831(.a(n12882), .b(n12881), .O(n12883));
  andx  g11832(.a(n12680), .b(n12883), .O(n12884));
  orx   g11833(.a(n12680), .b(n12883), .O(n12885));
  andx  g11834(.a(n12885), .b(n12675), .O(n12886));
  orx   g11835(.a(n12886), .b(n12884), .O(n12887));
  andx  g11836(.a(n12887), .b(n12880), .O(n12888));
  invx  g11837(.a(n12884), .O(n12889));
  andx  g11838(.a(n12685), .b(n12674), .O(n12890));
  orx   g11839(.a(n12890), .b(n12676), .O(n12891));
  andx  g11840(.a(n12891), .b(n12889), .O(n12892));
  andx  g11841(.a(n12892), .b(n12879), .O(n12893));
  orx   g11842(.a(n12893), .b(n12888), .O(n12894));
  andx  g11843(.a(n12894), .b(n12878), .O(n12895));
  orx   g11844(.a(n12894), .b(n12878), .O(n12896));
  invx  g11845(.a(n12896), .O(n12897));
  orx   g11846(.a(n12897), .b(n12895), .O(n12898));
  orx   g11847(.a(n12697), .b(n12691), .O(n12899));
  andx  g11848(.a(n12899), .b(n12702), .O(n12900));
  orx   g11849(.a(n12900), .b(n12000), .O(n12901));
  andx  g11850(.a(n12696), .b(n12701), .O(n12902));
  orx   g11851(.a(n12902), .b(n12694), .O(n12903));
  andx  g11852(.a(n11451), .b(n3180), .O(n12904));
  orx   g11853(.a(n12904), .b(n12903), .O(n12905));
  andx  g11854(.a(n12905), .b(n12901), .O(n12906));
  orx   g11855(.a(n12906), .b(n12898), .O(n12907));
  invx  g11856(.a(n12895), .O(n12908));
  andx  g11857(.a(n12896), .b(n12908), .O(n12909));
  andx  g11858(.a(n12903), .b(n11451), .O(n12910));
  invx  g11859(.a(n12904), .O(n12911));
  andx  g11860(.a(n12911), .b(n12900), .O(n12912));
  orx   g11861(.a(n12912), .b(n12910), .O(n12913));
  orx   g11862(.a(n12913), .b(n12909), .O(n12914));
  andx  g11863(.a(n12914), .b(n12907), .O(n12915));
  andx  g11864(.a(n12710), .b(n12722), .O(n12916));
  invx  g11865(.a(n12916), .O(n12917));
  orx   g11866(.a(n12715), .b(n12705), .O(n12918));
  andx  g11867(.a(n12918), .b(n12717), .O(n12919));
  andx  g11868(.a(n12919), .b(n12917), .O(n12920));
  orx   g11869(.a(n12920), .b(n12915), .O(n12921));
  andx  g11870(.a(n12913), .b(n12909), .O(n12922));
  andx  g11871(.a(n12906), .b(n12898), .O(n12923));
  orx   g11872(.a(n12923), .b(n12922), .O(n12924));
  andx  g11873(.a(n12709), .b(n12722), .O(n12925));
  orx   g11874(.a(n12925), .b(n12724), .O(n12926));
  orx   g11875(.a(n12926), .b(n12916), .O(n12927));
  orx   g11876(.a(n12927), .b(n12924), .O(n12928));
  andx  g11877(.a(n12928), .b(n12921), .O(n12929));
  andx  g11878(.a(n12737), .b(n12535), .O(n12930));
  andx  g11879(.a(n12727), .b(n12538), .O(n12931));
  orx   g11880(.a(n12931), .b(n12930), .O(n12932));
  andx  g11881(.a(n12742), .b(n12738), .O(n12933));
  orx   g11882(.a(n12933), .b(n12932), .O(n12934));
  andx  g11883(.a(n12934), .b(n12929), .O(n12935));
  andx  g11884(.a(n12927), .b(n12924), .O(n12936));
  andx  g11885(.a(n12920), .b(n12915), .O(n12937));
  orx   g11886(.a(n12937), .b(n12936), .O(n12938));
  invx  g11887(.a(n12934), .O(n12939));
  andx  g11888(.a(n12939), .b(n12938), .O(n12940));
  orx   g11889(.a(n12940), .b(n12935), .O(po15));
  invx  g11890(.a(n12931), .O(n12942));
  andx  g11891(.a(n12942), .b(n12734), .O(n12943));
  andx  g11892(.a(n12733), .b(n12536), .O(n12944));
  orx   g11893(.a(n12523), .b(n12520), .O(n12945));
  orx   g11894(.a(n12515), .b(n12306), .O(n12946));
  andx  g11895(.a(n12946), .b(n12945), .O(n12947));
  orx   g11896(.a(n12285), .b(n12044), .O(n12948));
  andx  g11897(.a(n12948), .b(n12947), .O(n12949));
  orx   g11898(.a(n12949), .b(n12042), .O(n12950));
  orx   g11899(.a(n12950), .b(n12292), .O(n12951));
  andx  g11900(.a(n12951), .b(n12529), .O(n12952));
  orx   g11901(.a(n12952), .b(n12944), .O(n12953));
  andx  g11902(.a(n12953), .b(n12943), .O(n12954));
  orx   g11903(.a(n12954), .b(n12929), .O(n12955));
  orx   g11904(.a(n12929), .b(n12944), .O(n12956));
  andx  g11905(.a(n12527), .b(n12287), .O(n12957));
  invx  g11906(.a(n12957), .O(n12958));
  orx   g11907(.a(n12958), .b(n12956), .O(n12959));
  orx   g11908(.a(n12959), .b(n12035), .O(n12960));
  andx  g11909(.a(n12960), .b(n12955), .O(n12961));
  orx   g11910(.a(n12920), .b(n12924), .O(n12962));
  orx   g11911(.a(n12912), .b(n12909), .O(n12963));
  andx  g11912(.a(n12963), .b(n12901), .O(n12964));
  andx  g11913(.a(n10356), .b(n3645), .O(n12965));
  andx  g11914(.a(n12829), .b(n12831), .O(n12966));
  orx   g11915(.a(n12966), .b(n12754), .O(n12967));
  orx   g11916(.a(n12967), .b(n12965), .O(n12968));
  orx   g11917(.a(n12836), .b(n12751), .O(n12969));
  andx  g11918(.a(n12969), .b(n12832), .O(n12970));
  orx   g11919(.a(n12970), .b(n11053), .O(n12971));
  andx  g11920(.a(n12971), .b(n12968), .O(n12972));
  andx  g11921(.a(n9470), .b(n4063), .O(n12973));
  andx  g11922(.a(n12805), .b(n12759), .O(n12974));
  orx   g11923(.a(n12974), .b(n12801), .O(n12975));
  orx   g11924(.a(n12975), .b(n12973), .O(n12976));
  invx  g11925(.a(n12976), .O(n12977));
  andx  g11926(.a(n12975), .b(n9470), .O(n12978));
  orx   g11927(.a(n12978), .b(n12977), .O(n12979));
  andx  g11928(.a(n11157), .b(n8852), .O(n12987));
  invx  g11929(.a(n12987), .O(n12988));
  andx  g11930(.a(n12988), .b(n12769), .O(n12989));
  orx   g11931(.a(n12989), .b(n10161), .O(n12990));
  andx  g11932(.a(n12768), .b(n8852), .O(n12991));
  invx  g11933(.a(n12991), .O(n12992));
  andx  g11934(.a(n12992), .b(n12990), .O(n12993));
  andx  g11935(.a(n9267), .b(n4114), .O(n12999));
  andx  g11936(.a(n12788), .b(n11260), .O(n13003));
  orx   g11937(.a(n13003), .b(n12783), .O(n13004));
  andx  g11938(.a(n13004), .b(n12787), .O(n13005));
  invx  g11939(.a(n13005), .O(n13006));
  andx  g11940(.a(n13006), .b(n12999), .O(n13007));
  invx  g11941(.a(n12999), .O(n13008));
  andx  g11942(.a(n13005), .b(n13008), .O(n13009));
  orx   g11943(.a(n13009), .b(n13007), .O(n13010));
  orx   g11944(.a(n13010), .b(n9050), .O(n13011));
  invx  g11945(.a(n13011), .O(n13012));
  andx  g11946(.a(n13010), .b(n9050), .O(n13013));
  orx   g11947(.a(n13013), .b(n13012), .O(n13014));
  andx  g11948(.a(n13014), .b(n12979), .O(n13015));
  invx  g11949(.a(n12978), .O(n13016));
  andx  g11950(.a(n13016), .b(n12976), .O(n13017));
  invx  g11951(.a(n13013), .O(n13018));
  andx  g11952(.a(n13018), .b(n13011), .O(n13019));
  andx  g11953(.a(n13019), .b(n13017), .O(n13020));
  orx   g11954(.a(n13020), .b(n13015), .O(n13021));
  andx  g11955(.a(n12811), .b(n12824), .O(n13022));
  invx  g11956(.a(n13022), .O(n13023));
  andx  g11957(.a(n12817), .b(n12807), .O(n13024));
  orx   g11958(.a(n13024), .b(n12818), .O(n13025));
  andx  g11959(.a(n13025), .b(n13023), .O(n13026));
  andx  g11960(.a(n7902), .b(n3721), .O(n13027));
  invx  g11961(.a(n13027), .O(n13028));
  andx  g11962(.a(n13028), .b(n13026), .O(n13029));
  orx   g11963(.a(n12811), .b(n12824), .O(n13030));
  andx  g11964(.a(n13030), .b(n12812), .O(n13031));
  orx   g11965(.a(n13031), .b(n13022), .O(n13032));
  andx  g11966(.a(n13027), .b(n13032), .O(n13033));
  orx   g11967(.a(n13033), .b(n13029), .O(n13034));
  orx   g11968(.a(n13034), .b(n13021), .O(n13035));
  orx   g11969(.a(n13019), .b(n13017), .O(n13036));
  orx   g11970(.a(n13014), .b(n12979), .O(n13037));
  andx  g11971(.a(n13037), .b(n13036), .O(n13038));
  orx   g11972(.a(n13027), .b(n13032), .O(n13039));
  orx   g11973(.a(n13028), .b(n13026), .O(n13040));
  andx  g11974(.a(n13040), .b(n13039), .O(n13041));
  orx   g11975(.a(n13041), .b(n13038), .O(n13042));
  andx  g11976(.a(n13042), .b(n13035), .O(n13043));
  orx   g11977(.a(n13043), .b(n12972), .O(n13044));
  invx  g11978(.a(n12965), .O(n13045));
  andx  g11979(.a(n12970), .b(n13045), .O(n13046));
  andx  g11980(.a(n12967), .b(n10356), .O(n13047));
  orx   g11981(.a(n13047), .b(n13046), .O(n13048));
  andx  g11982(.a(n13041), .b(n13038), .O(n13049));
  andx  g11983(.a(n13034), .b(n13021), .O(n13050));
  orx   g11984(.a(n13050), .b(n13049), .O(n13051));
  orx   g11985(.a(n13051), .b(n13048), .O(n13052));
  andx  g11986(.a(n13052), .b(n13044), .O(n13053));
  andx  g11987(.a(n10751), .b(n3413), .O(n13054));
  invx  g11988(.a(n13054), .O(n13055));
  andx  g11989(.a(n12849), .b(n12838), .O(n13056));
  orx   g11990(.a(n12849), .b(n12838), .O(n13057));
  andx  g11991(.a(n13057), .b(n12839), .O(n13058));
  orx   g11992(.a(n13058), .b(n13056), .O(n13059));
  andx  g11993(.a(n13059), .b(n13055), .O(n13060));
  invx  g11994(.a(n13056), .O(n13061));
  andx  g11995(.a(n12844), .b(n12855), .O(n13062));
  orx   g11996(.a(n13062), .b(n12846), .O(n13063));
  andx  g11997(.a(n13063), .b(n13061), .O(n13064));
  andx  g11998(.a(n13064), .b(n13054), .O(n13065));
  orx   g11999(.a(n13065), .b(n13060), .O(n13066));
  andx  g12000(.a(n13066), .b(n13053), .O(n13067));
  andx  g12001(.a(n13051), .b(n13048), .O(n13068));
  andx  g12002(.a(n13043), .b(n12972), .O(n13069));
  orx   g12003(.a(n13069), .b(n13068), .O(n13070));
  orx   g12004(.a(n13064), .b(n13054), .O(n13071));
  orx   g12005(.a(n13059), .b(n13055), .O(n13072));
  andx  g12006(.a(n13072), .b(n13071), .O(n13073));
  andx  g12007(.a(n13073), .b(n13070), .O(n13074));
  orx   g12008(.a(n13074), .b(n13067), .O(n13075));
  orx   g12009(.a(n12868), .b(n12860), .O(n13076));
  andx  g12010(.a(n13076), .b(n12874), .O(n13077));
  orx   g12011(.a(n13077), .b(n11714), .O(n13078));
  andx  g12012(.a(n12875), .b(n12873), .O(n13079));
  orx   g12013(.a(n13079), .b(n12863), .O(n13080));
  andx  g12014(.a(n11120), .b(n3171), .O(n13081));
  orx   g12015(.a(n13081), .b(n13080), .O(n13082));
  andx  g12016(.a(n13082), .b(n13078), .O(n13083));
  orx   g12017(.a(n13083), .b(n13075), .O(n13084));
  orx   g12018(.a(n13073), .b(n13070), .O(n13085));
  orx   g12019(.a(n13066), .b(n13053), .O(n13086));
  andx  g12020(.a(n13086), .b(n13085), .O(n13087));
  andx  g12021(.a(n13080), .b(n11120), .O(n13088));
  invx  g12022(.a(n13081), .O(n13089));
  andx  g12023(.a(n13089), .b(n13077), .O(n13090));
  orx   g12024(.a(n13090), .b(n13088), .O(n13091));
  orx   g12025(.a(n13091), .b(n13087), .O(n13092));
  andx  g12026(.a(n13092), .b(n13084), .O(n13093));
  andx  g12027(.a(n11451), .b(n3429), .O(n13094));
  invx  g12028(.a(n13094), .O(n13095));
  orx   g12029(.a(n12876), .b(n12873), .O(n13096));
  orx   g12030(.a(n12869), .b(n12860), .O(n13097));
  andx  g12031(.a(n13097), .b(n13096), .O(n13098));
  andx  g12032(.a(n12887), .b(n13098), .O(n13099));
  invx  g12033(.a(n13099), .O(n13100));
  andx  g12034(.a(n12892), .b(n12878), .O(n13101));
  orx   g12035(.a(n13101), .b(n12880), .O(n13102));
  andx  g12036(.a(n13102), .b(n13100), .O(n13103));
  orx   g12037(.a(n13103), .b(n13095), .O(n13104));
  orx   g12038(.a(n12887), .b(n13098), .O(n13105));
  andx  g12039(.a(n13105), .b(n12879), .O(n13106));
  orx   g12040(.a(n13106), .b(n13099), .O(n13107));
  orx   g12041(.a(n13107), .b(n13094), .O(n13108));
  andx  g12042(.a(n13108), .b(n13104), .O(n13109));
  andx  g12043(.a(n13109), .b(n13093), .O(n13110));
  andx  g12044(.a(n13091), .b(n13087), .O(n13111));
  andx  g12045(.a(n13083), .b(n13075), .O(n13112));
  orx   g12046(.a(n13112), .b(n13111), .O(n13113));
  andx  g12047(.a(n13107), .b(n13094), .O(n13114));
  andx  g12048(.a(n13103), .b(n13095), .O(n13115));
  orx   g12049(.a(n13115), .b(n13114), .O(n13116));
  andx  g12050(.a(n13116), .b(n13113), .O(n13117));
  orx   g12051(.a(n13117), .b(n13110), .O(n13118));
  andx  g12052(.a(n13118), .b(n12964), .O(n13119));
  andx  g12053(.a(n12905), .b(n12898), .O(n13120));
  orx   g12054(.a(n13120), .b(n12910), .O(n13121));
  orx   g12055(.a(n13116), .b(n13113), .O(n13122));
  orx   g12056(.a(n13109), .b(n13093), .O(n13123));
  andx  g12057(.a(n13123), .b(n13122), .O(n13124));
  andx  g12058(.a(n13124), .b(n13121), .O(n13125));
  orx   g12059(.a(n13125), .b(n13119), .O(n13126));
  invx  g12060(.a(n13126), .O(n13127));
  andx  g12061(.a(n13127), .b(n12962), .O(n13128));
  andx  g12062(.a(n13128), .b(n12961), .O(n13129));
  andx  g12063(.a(n12927), .b(n12915), .O(n13130));
  andx  g12064(.a(n13126), .b(n13130), .O(n13131));
  andx  g12065(.a(n12527), .b(n12023), .O(n13132));
  andx  g12066(.a(n13132), .b(n12287), .O(n13133));
  orx   g12067(.a(n13133), .b(n12528), .O(n13134));
  andx  g12068(.a(n13134), .b(n12738), .O(n13135));
  orx   g12069(.a(n13135), .b(n12932), .O(n13136));
  andx  g12070(.a(n13136), .b(n12938), .O(n13137));
  andx  g12071(.a(n12938), .b(n12738), .O(n13138));
  andx  g12072(.a(n12957), .b(n13138), .O(n13139));
  andx  g12073(.a(n13139), .b(n12296), .O(n13140));
  orx   g12074(.a(n13140), .b(n13137), .O(n13141));
  andx  g12075(.a(n13126), .b(n13141), .O(n13142));
  orx   g12076(.a(n13142), .b(n13131), .O(n13143));
  orx   g12077(.a(n13143), .b(n13129), .O(po16));
  andx  g12078(.a(n10751), .b(n3645), .O(n13145));
  andx  g12079(.a(n13051), .b(n12968), .O(n13146));
  orx   g12080(.a(n13146), .b(n13047), .O(n13147));
  orx   g12081(.a(n13147), .b(n13145), .O(n13148));
  andx  g12082(.a(n13147), .b(n10751), .O(n13149));
  invx  g12083(.a(n13149), .O(n13150));
  andx  g12084(.a(n13150), .b(n13148), .O(n13151));
  andx  g12085(.a(n7902), .b(n4063), .O(n13152));
  invx  g12086(.a(n13152), .O(n13153));
  orx   g12087(.a(n13019), .b(n12977), .O(n13154));
  andx  g12088(.a(n13154), .b(n13016), .O(n13155));
  andx  g12089(.a(n13155), .b(n13153), .O(n13156));
  andx  g12090(.a(n13014), .b(n12976), .O(n13157));
  orx   g12091(.a(n13157), .b(n12978), .O(n13158));
  andx  g12092(.a(n13158), .b(n7902), .O(n13159));
  orx   g12093(.a(n13159), .b(n13156), .O(n13160));
  andx  g12094(.a(n12993), .b(n12988), .O(n13161));
  orx   g12095(.a(n13161), .b(n10585), .O(n13162));
  orx   g12096(.a(n12993), .b(n11260), .O(n13163));
  andx  g12097(.a(n13163), .b(n13162), .O(n13164));
  andx  g12098(.a(n9470), .b(n4114), .O(n13176));
  invx  g12099(.a(n13176), .O(n13177));
  andx  g12100(.a(n13006), .b(n9050), .O(n13178));
  invx  g12101(.a(n13178), .O(n13179));
  andx  g12102(.a(n13005), .b(n10585), .O(n13180));
  orx   g12103(.a(n13180), .b(n13008), .O(n13181));
  andx  g12104(.a(n13181), .b(n13179), .O(n13182));
  orx   g12105(.a(n13182), .b(n13177), .O(n13183));
  andx  g12106(.a(n13182), .b(n13177), .O(n13184));
  invx  g12107(.a(n13184), .O(n13185));
  andx  g12108(.a(n13185), .b(n13183), .O(n13186));
  andx  g12109(.a(n13186), .b(n9266), .O(n13187));
  invx  g12110(.a(n13183), .O(n13189));
  orx   g12111(.a(n13184), .b(n13189), .O(n13190));
  andx  g12112(.a(n13190), .b(n9267), .O(n13191));
  orx   g12113(.a(n13191), .b(n13187), .O(n13192));
  andx  g12114(.a(n13192), .b(n13160), .O(n13193));
  orx   g12115(.a(n13158), .b(n13152), .O(n13194));
  orx   g12116(.a(n13155), .b(n11349), .O(n13195));
  andx  g12117(.a(n13195), .b(n13194), .O(n13196));
  orx   g12118(.a(n13190), .b(n9267), .O(n13197));
  orx   g12119(.a(n13186), .b(n9266), .O(n13198));
  andx  g12120(.a(n13198), .b(n13197), .O(n13199));
  andx  g12121(.a(n13199), .b(n13196), .O(n13200));
  orx   g12122(.a(n13200), .b(n13193), .O(n13201));
  andx  g12123(.a(n13032), .b(n13021), .O(n13202));
  invx  g12124(.a(n13202), .O(n13203));
  andx  g12125(.a(n13026), .b(n13038), .O(n13204));
  orx   g12126(.a(n13204), .b(n13028), .O(n13205));
  andx  g12127(.a(n13205), .b(n13203), .O(n13206));
  andx  g12128(.a(n10356), .b(n3721), .O(n13207));
  invx  g12129(.a(n13207), .O(n13208));
  andx  g12130(.a(n13208), .b(n13206), .O(n13209));
  orx   g12131(.a(n13032), .b(n13021), .O(n13210));
  andx  g12132(.a(n13210), .b(n13027), .O(n13211));
  orx   g12133(.a(n13211), .b(n13202), .O(n13212));
  andx  g12134(.a(n13207), .b(n13212), .O(n13213));
  orx   g12135(.a(n13213), .b(n13209), .O(n13214));
  orx   g12136(.a(n13214), .b(n13201), .O(n13215));
  orx   g12137(.a(n13199), .b(n13196), .O(n13216));
  orx   g12138(.a(n13192), .b(n13160), .O(n13217));
  andx  g12139(.a(n13217), .b(n13216), .O(n13218));
  orx   g12140(.a(n13207), .b(n13212), .O(n13219));
  orx   g12141(.a(n13208), .b(n13206), .O(n13220));
  andx  g12142(.a(n13220), .b(n13219), .O(n13221));
  orx   g12143(.a(n13221), .b(n13218), .O(n13222));
  andx  g12144(.a(n13222), .b(n13215), .O(n13223));
  orx   g12145(.a(n13223), .b(n13151), .O(n13224));
  invx  g12146(.a(n13148), .O(n13225));
  orx   g12147(.a(n13149), .b(n13225), .O(n13226));
  andx  g12148(.a(n13221), .b(n13218), .O(n13227));
  andx  g12149(.a(n13214), .b(n13201), .O(n13228));
  orx   g12150(.a(n13228), .b(n13227), .O(n13229));
  orx   g12151(.a(n13229), .b(n13226), .O(n13230));
  andx  g12152(.a(n13230), .b(n13224), .O(n13231));
  andx  g12153(.a(n11120), .b(n3413), .O(n13232));
  invx  g12154(.a(n13232), .O(n13233));
  andx  g12155(.a(n13059), .b(n13070), .O(n13234));
  orx   g12156(.a(n13059), .b(n13070), .O(n13235));
  andx  g12157(.a(n13235), .b(n13054), .O(n13236));
  orx   g12158(.a(n13236), .b(n13234), .O(n13237));
  andx  g12159(.a(n13237), .b(n13233), .O(n13238));
  invx  g12160(.a(n13234), .O(n13239));
  andx  g12161(.a(n13064), .b(n13053), .O(n13240));
  orx   g12162(.a(n13240), .b(n13055), .O(n13241));
  andx  g12163(.a(n13241), .b(n13239), .O(n13242));
  andx  g12164(.a(n13242), .b(n13232), .O(n13243));
  orx   g12165(.a(n13243), .b(n13238), .O(n13244));
  andx  g12166(.a(n13244), .b(n13231), .O(n13245));
  andx  g12167(.a(n13229), .b(n13226), .O(n13246));
  andx  g12168(.a(n13223), .b(n13151), .O(n13247));
  orx   g12169(.a(n13247), .b(n13246), .O(n13248));
  orx   g12170(.a(n13242), .b(n13232), .O(n13249));
  orx   g12171(.a(n13237), .b(n13233), .O(n13250));
  andx  g12172(.a(n13250), .b(n13249), .O(n13251));
  andx  g12173(.a(n13251), .b(n13248), .O(n13252));
  orx   g12174(.a(n13252), .b(n13245), .O(n13253));
  orx   g12175(.a(n13090), .b(n13087), .O(n13254));
  andx  g12176(.a(n13254), .b(n13078), .O(n13255));
  orx   g12177(.a(n13255), .b(n12000), .O(n13256));
  andx  g12178(.a(n13082), .b(n13075), .O(n13257));
  orx   g12179(.a(n13257), .b(n13088), .O(n13258));
  andx  g12180(.a(n11451), .b(n3171), .O(n13259));
  orx   g12181(.a(n13259), .b(n13258), .O(n13260));
  andx  g12182(.a(n13260), .b(n13256), .O(n13261));
  orx   g12183(.a(n13261), .b(n13253), .O(n13262));
  orx   g12184(.a(n13251), .b(n13248), .O(n13263));
  orx   g12185(.a(n13244), .b(n13231), .O(n13264));
  andx  g12186(.a(n13264), .b(n13263), .O(n13265));
  andx  g12187(.a(n13258), .b(n11451), .O(n13266));
  invx  g12188(.a(n13259), .O(n13267));
  andx  g12189(.a(n13267), .b(n13255), .O(n13268));
  orx   g12190(.a(n13268), .b(n13266), .O(n13269));
  orx   g12191(.a(n13269), .b(n13265), .O(n13270));
  andx  g12192(.a(n13270), .b(n13262), .O(n13271));
  andx  g12193(.a(n13094), .b(n13093), .O(n13272));
  invx  g12194(.a(n13272), .O(n13273));
  andx  g12195(.a(n13095), .b(n13113), .O(n13274));
  orx   g12196(.a(n13274), .b(n13103), .O(n13275));
  andx  g12197(.a(n13275), .b(n13273), .O(n13276));
  andx  g12198(.a(n13276), .b(n13271), .O(n13277));
  andx  g12199(.a(n13269), .b(n13265), .O(n13278));
  andx  g12200(.a(n13261), .b(n13253), .O(n13279));
  orx   g12201(.a(n13279), .b(n13278), .O(n13280));
  orx   g12202(.a(n13094), .b(n13093), .O(n13281));
  andx  g12203(.a(n13281), .b(n13107), .O(n13282));
  orx   g12204(.a(n13282), .b(n13272), .O(n13283));
  andx  g12205(.a(n13283), .b(n13280), .O(n13284));
  orx   g12206(.a(n13284), .b(n13277), .O(n13285));
  orx   g12207(.a(n13285), .b(n13125), .O(n13286));
  andx  g12208(.a(n13285), .b(n13125), .O(n13287));
  invx  g12209(.a(n13287), .O(n13288));
  andx  g12210(.a(n13288), .b(n13286), .O(n13289));
  invx  g12211(.a(n13289), .O(n13290));
  andx  g12212(.a(n12962), .b(n12961), .O(n13291));
  orx   g12213(.a(n13291), .b(n13126), .O(n13292));
  orx   g12214(.a(n13292), .b(n13290), .O(n13293));
  invx  g12215(.a(n13292), .O(n13294));
  orx   g12216(.a(n13294), .b(n13289), .O(n13295));
  andx  g12217(.a(n13295), .b(n13293), .O(po17));
  andx  g12218(.a(n13283), .b(n13271), .O(n13297));
  invx  g12219(.a(n13297), .O(n13298));
  andx  g12220(.a(n13260), .b(n13253), .O(n13299));
  orx   g12221(.a(n13299), .b(n13266), .O(n13300));
  invx  g12222(.a(n13300), .O(n13301));
  andx  g12223(.a(n11120), .b(n3645), .O(n13302));
  andx  g12224(.a(n13229), .b(n13148), .O(n13303));
  orx   g12225(.a(n13303), .b(n13149), .O(n13304));
  orx   g12226(.a(n13304), .b(n13302), .O(n13305));
  invx  g12227(.a(n13305), .O(n13306));
  andx  g12228(.a(n13304), .b(n11120), .O(n13307));
  orx   g12229(.a(n13307), .b(n13306), .O(n13308));
  andx  g12230(.a(n10356), .b(n4063), .O(n13309));
  invx  g12231(.a(n13309), .O(n13310));
  orx   g12232(.a(n13199), .b(n13156), .O(n13311));
  andx  g12233(.a(n13311), .b(n13195), .O(n13312));
  andx  g12234(.a(n13312), .b(n13310), .O(n13313));
  andx  g12235(.a(n13192), .b(n13194), .O(n13314));
  orx   g12236(.a(n13314), .b(n13159), .O(n13315));
  andx  g12237(.a(n13315), .b(n10356), .O(n13316));
  orx   g12238(.a(n13316), .b(n13313), .O(n13317));
  andx  g12239(.a(n2429), .b(n9470), .O(n13320));
  andx  g12240(.a(n2724), .b(n9267), .O(n13323));
  orx   g12241(.a(n13323), .b(n13320), .O(n13324));
  invx  g12242(.a(n13164), .O(n13325));
  andx  g12243(.a(n11157), .b(n9267), .O(n13326));
  orx   g12244(.a(n13326), .b(n13325), .O(n13327));
  andx  g12245(.a(n13327), .b(n9050), .O(n13328));
  andx  g12246(.a(n13325), .b(n9267), .O(n13329));
  orx   g12247(.a(n13329), .b(n13328), .O(n13330));
  invx  g12248(.a(n13330), .O(n13331));
  andx  g12249(.a(n13331), .b(n13324), .O(n13332));
  invx  g12250(.a(n13332), .O(n13333));
  orx   g12251(.a(n13331), .b(n13324), .O(n13334));
  andx  g12252(.a(n13334), .b(n13333), .O(n13335));
  invx  g12253(.a(n13182), .O(n13336));
  andx  g12254(.a(n13336), .b(n9267), .O(n13337));
  andx  g12255(.a(n13182), .b(n9266), .O(n13338));
  orx   g12256(.a(n13338), .b(n13177), .O(n13339));
  invx  g12257(.a(n13339), .O(n13340));
  orx   g12258(.a(n13340), .b(n13337), .O(n13341));
  andx  g12259(.a(n7902), .b(n4114), .O(n13342));
  orx   g12260(.a(n13342), .b(n13341), .O(n13343));
  invx  g12261(.a(n13337), .O(n13344));
  andx  g12262(.a(n13339), .b(n13344), .O(n13345));
  invx  g12263(.a(n13342), .O(n13346));
  orx   g12264(.a(n13346), .b(n13345), .O(n13347));
  andx  g12265(.a(n13347), .b(n13343), .O(n13348));
  andx  g12266(.a(n13348), .b(n13335), .O(n13349));
  invx  g12267(.a(n13335), .O(n13350));
  andx  g12268(.a(n13346), .b(n13345), .O(n13351));
  andx  g12269(.a(n13342), .b(n13341), .O(n13352));
  orx   g12270(.a(n13352), .b(n13351), .O(n13353));
  andx  g12271(.a(n13353), .b(n13350), .O(n13354));
  orx   g12272(.a(n13354), .b(n13349), .O(n13355));
  andx  g12273(.a(n13355), .b(n13317), .O(n13356));
  orx   g12274(.a(n13315), .b(n13309), .O(n13357));
  orx   g12275(.a(n13312), .b(n11053), .O(n13358));
  andx  g12276(.a(n13358), .b(n13357), .O(n13359));
  orx   g12277(.a(n13353), .b(n13350), .O(n13360));
  orx   g12278(.a(n13348), .b(n13335), .O(n13361));
  andx  g12279(.a(n13361), .b(n13360), .O(n13362));
  andx  g12280(.a(n13362), .b(n13359), .O(n13363));
  orx   g12281(.a(n13363), .b(n13356), .O(n13364));
  andx  g12282(.a(n13212), .b(n13201), .O(n13365));
  invx  g12283(.a(n13365), .O(n13366));
  andx  g12284(.a(n13206), .b(n13218), .O(n13367));
  orx   g12285(.a(n13367), .b(n13208), .O(n13368));
  andx  g12286(.a(n13368), .b(n13366), .O(n13369));
  andx  g12287(.a(n10751), .b(n3721), .O(n13370));
  invx  g12288(.a(n13370), .O(n13371));
  andx  g12289(.a(n13371), .b(n13369), .O(n13372));
  orx   g12290(.a(n13212), .b(n13201), .O(n13373));
  andx  g12291(.a(n13373), .b(n13207), .O(n13374));
  orx   g12292(.a(n13374), .b(n13365), .O(n13375));
  andx  g12293(.a(n13370), .b(n13375), .O(n13376));
  orx   g12294(.a(n13376), .b(n13372), .O(n13377));
  orx   g12295(.a(n13377), .b(n13364), .O(n13378));
  orx   g12296(.a(n13362), .b(n13359), .O(n13379));
  orx   g12297(.a(n13355), .b(n13317), .O(n13380));
  andx  g12298(.a(n13380), .b(n13379), .O(n13381));
  orx   g12299(.a(n13370), .b(n13375), .O(n13382));
  orx   g12300(.a(n13371), .b(n13369), .O(n13383));
  andx  g12301(.a(n13383), .b(n13382), .O(n13384));
  orx   g12302(.a(n13384), .b(n13381), .O(n13385));
  andx  g12303(.a(n13385), .b(n13378), .O(n13386));
  andx  g12304(.a(n13386), .b(n13308), .O(n13387));
  invx  g12305(.a(n13307), .O(n13388));
  andx  g12306(.a(n13388), .b(n13305), .O(n13389));
  andx  g12307(.a(n13384), .b(n13381), .O(n13390));
  andx  g12308(.a(n13377), .b(n13364), .O(n13391));
  orx   g12309(.a(n13391), .b(n13390), .O(n13392));
  andx  g12310(.a(n13392), .b(n13389), .O(n13393));
  orx   g12311(.a(n13393), .b(n13387), .O(n13394));
  andx  g12312(.a(n11451), .b(n3413), .O(n13395));
  invx  g12313(.a(n13395), .O(n13396));
  andx  g12314(.a(n13237), .b(n13248), .O(n13397));
  orx   g12315(.a(n13237), .b(n13248), .O(n13398));
  andx  g12316(.a(n13398), .b(n13232), .O(n13399));
  orx   g12317(.a(n13399), .b(n13397), .O(n13400));
  andx  g12318(.a(n13400), .b(n13396), .O(n13401));
  invx  g12319(.a(n13397), .O(n13402));
  andx  g12320(.a(n13242), .b(n13231), .O(n13403));
  orx   g12321(.a(n13403), .b(n13233), .O(n13404));
  andx  g12322(.a(n13404), .b(n13402), .O(n13405));
  andx  g12323(.a(n13405), .b(n13395), .O(n13406));
  orx   g12324(.a(n13406), .b(n13401), .O(n13407));
  andx  g12325(.a(n13407), .b(n13394), .O(n13408));
  orx   g12326(.a(n13392), .b(n13389), .O(n13409));
  orx   g12327(.a(n13386), .b(n13308), .O(n13410));
  andx  g12328(.a(n13410), .b(n13409), .O(n13411));
  orx   g12329(.a(n13405), .b(n13395), .O(n13412));
  orx   g12330(.a(n13400), .b(n13396), .O(n13413));
  andx  g12331(.a(n13413), .b(n13412), .O(n13414));
  andx  g12332(.a(n13414), .b(n13411), .O(n13415));
  orx   g12333(.a(n13415), .b(n13408), .O(n13416));
  orx   g12334(.a(n13416), .b(n13301), .O(n13417));
  orx   g12335(.a(n13414), .b(n13411), .O(n13418));
  orx   g12336(.a(n13407), .b(n13394), .O(n13419));
  andx  g12337(.a(n13419), .b(n13418), .O(n13420));
  orx   g12338(.a(n13420), .b(n13300), .O(n13421));
  andx  g12339(.a(n13421), .b(n13417), .O(n13422));
  orx   g12340(.a(n13422), .b(n13298), .O(n13423));
  andx  g12341(.a(n13420), .b(n13300), .O(n13424));
  andx  g12342(.a(n13416), .b(n13301), .O(n13425));
  orx   g12343(.a(n13425), .b(n13424), .O(n13426));
  orx   g12344(.a(n13426), .b(n13297), .O(n13427));
  andx  g12345(.a(n13427), .b(n13423), .O(n13428));
  invx  g12346(.a(n13428), .O(n13429));
  orx   g12347(.a(n13118), .b(n12964), .O(n13430));
  orx   g12348(.a(n13283), .b(n13280), .O(n13431));
  orx   g12349(.a(n13276), .b(n13271), .O(n13432));
  andx  g12350(.a(n13432), .b(n13431), .O(n13433));
  andx  g12351(.a(n13433), .b(n13430), .O(n13434));
  andx  g12352(.a(n13293), .b(n13288), .O(n13436));
  invx  g12353(.a(n13436), .O(n13437));
  andx  g12354(.a(n13437), .b(n13429), .O(n13438));
  andx  g12355(.a(n13436), .b(n13428), .O(n13439));
  orx   g12356(.a(n13439), .b(n13438), .O(po18));
  andx  g12357(.a(n13395), .b(n13411), .O(n13441));
  andx  g12358(.a(n13400), .b(n13411), .O(n13442));
  andx  g12359(.a(n13400), .b(n13395), .O(n13443));
  orx   g12360(.a(n13443), .b(n13442), .O(n13444));
  orx   g12361(.a(n13444), .b(n13441), .O(n13445));
  andx  g12362(.a(n11451), .b(n3645), .O(n13446));
  andx  g12363(.a(n13392), .b(n13305), .O(n13447));
  orx   g12364(.a(n13447), .b(n13307), .O(n13448));
  orx   g12365(.a(n13448), .b(n13446), .O(n13449));
  orx   g12366(.a(n13386), .b(n13306), .O(n13450));
  andx  g12367(.a(n13450), .b(n13388), .O(n13451));
  orx   g12368(.a(n13451), .b(n12000), .O(n13452));
  andx  g12369(.a(n13452), .b(n13449), .O(n13453));
  andx  g12370(.a(n10751), .b(n4063), .O(n13454));
  invx  g12371(.a(n13454), .O(n13455));
  orx   g12372(.a(n13362), .b(n13313), .O(n13456));
  andx  g12373(.a(n13456), .b(n13358), .O(n13457));
  andx  g12374(.a(n13457), .b(n13455), .O(n13458));
  andx  g12375(.a(n13355), .b(n13357), .O(n13459));
  orx   g12376(.a(n13459), .b(n13316), .O(n13460));
  andx  g12377(.a(n13460), .b(n10751), .O(n13461));
  orx   g12378(.a(n13461), .b(n13458), .O(n13462));
  andx  g12379(.a(n11157), .b(n9470), .O(n13463));
  orx   g12380(.a(n13463), .b(n13330), .O(n13464));
  andx  g12381(.a(n13464), .b(n9267), .O(n13465));
  andx  g12382(.a(n13330), .b(n9470), .O(n13466));
  orx   g12383(.a(n13466), .b(n13465), .O(n13467));
  invx  g12384(.a(n13467), .O(n13468));
  andx  g12385(.a(n2724), .b(n9470), .O(n13471));
  andx  g12386(.a(n2429), .b(n7902), .O(n13474));
  orx   g12387(.a(n13474), .b(n13471), .O(n13475));
  andx  g12388(.a(n13475), .b(n13468), .O(n13476));
  invx  g12389(.a(n13476), .O(n13477));
  orx   g12390(.a(n13475), .b(n13468), .O(n13478));
  andx  g12391(.a(n13478), .b(n13477), .O(n13479));
  andx  g12392(.a(n13341), .b(n13350), .O(n13480));
  orx   g12393(.a(n13341), .b(n13350), .O(n13481));
  andx  g12394(.a(n13481), .b(n13342), .O(n13482));
  orx   g12395(.a(n13482), .b(n13480), .O(n13483));
  andx  g12396(.a(n10356), .b(n4114), .O(n13484));
  orx   g12397(.a(n13484), .b(n13483), .O(n13485));
  invx  g12398(.a(n13480), .O(n13486));
  andx  g12399(.a(n13345), .b(n13335), .O(n13487));
  orx   g12400(.a(n13487), .b(n13346), .O(n13488));
  andx  g12401(.a(n13488), .b(n13486), .O(n13489));
  invx  g12402(.a(n13484), .O(n13490));
  orx   g12403(.a(n13490), .b(n13489), .O(n13491));
  andx  g12404(.a(n13491), .b(n13485), .O(n13492));
  andx  g12405(.a(n13492), .b(n13479), .O(n13493));
  invx  g12406(.a(n13479), .O(n13494));
  andx  g12407(.a(n13490), .b(n13489), .O(n13495));
  andx  g12408(.a(n13484), .b(n13483), .O(n13496));
  orx   g12409(.a(n13496), .b(n13495), .O(n13497));
  andx  g12410(.a(n13497), .b(n13494), .O(n13498));
  orx   g12411(.a(n13498), .b(n13493), .O(n13499));
  andx  g12412(.a(n13499), .b(n13462), .O(n13500));
  orx   g12413(.a(n13460), .b(n13454), .O(n13501));
  orx   g12414(.a(n13457), .b(n11380), .O(n13502));
  andx  g12415(.a(n13502), .b(n13501), .O(n13503));
  orx   g12416(.a(n13497), .b(n13494), .O(n13504));
  orx   g12417(.a(n13492), .b(n13479), .O(n13505));
  andx  g12418(.a(n13505), .b(n13504), .O(n13506));
  andx  g12419(.a(n13506), .b(n13503), .O(n13507));
  orx   g12420(.a(n13507), .b(n13500), .O(n13508));
  andx  g12421(.a(n13375), .b(n13364), .O(n13509));
  invx  g12422(.a(n13509), .O(n13510));
  andx  g12423(.a(n13369), .b(n13381), .O(n13511));
  orx   g12424(.a(n13511), .b(n13371), .O(n13512));
  andx  g12425(.a(n13512), .b(n13510), .O(n13513));
  andx  g12426(.a(n11120), .b(n3721), .O(n13514));
  invx  g12427(.a(n13514), .O(n13515));
  andx  g12428(.a(n13515), .b(n13513), .O(n13516));
  orx   g12429(.a(n13375), .b(n13364), .O(n13517));
  andx  g12430(.a(n13517), .b(n13370), .O(n13518));
  orx   g12431(.a(n13518), .b(n13509), .O(n13519));
  andx  g12432(.a(n13514), .b(n13519), .O(n13520));
  orx   g12433(.a(n13520), .b(n13516), .O(n13521));
  orx   g12434(.a(n13521), .b(n13508), .O(n13522));
  andx  g12435(.a(n13521), .b(n13508), .O(n13523));
  invx  g12436(.a(n13523), .O(n13524));
  andx  g12437(.a(n13524), .b(n13522), .O(n13525));
  orx   g12438(.a(n13525), .b(n13453), .O(n13526));
  invx  g12439(.a(n13446), .O(n13527));
  andx  g12440(.a(n13451), .b(n13527), .O(n13528));
  andx  g12441(.a(n13448), .b(n11451), .O(n13529));
  orx   g12442(.a(n13529), .b(n13528), .O(n13530));
  invx  g12443(.a(n13522), .O(n13531));
  orx   g12444(.a(n13523), .b(n13531), .O(n13532));
  orx   g12445(.a(n13532), .b(n13530), .O(n13533));
  andx  g12446(.a(n13533), .b(n13526), .O(n13534));
  orx   g12447(.a(n13534), .b(n13445), .O(n13535));
  invx  g12448(.a(n13441), .O(n13536));
  orx   g12449(.a(n13405), .b(n13394), .O(n13537));
  invx  g12450(.a(n13443), .O(n13538));
  andx  g12451(.a(n13538), .b(n13537), .O(n13539));
  andx  g12452(.a(n13539), .b(n13536), .O(n13540));
  andx  g12453(.a(n13532), .b(n13530), .O(n13541));
  andx  g12454(.a(n13525), .b(n13453), .O(n13542));
  orx   g12455(.a(n13542), .b(n13541), .O(n13543));
  orx   g12456(.a(n13543), .b(n13540), .O(n13544));
  andx  g12457(.a(n13544), .b(n13535), .O(n13545));
  andx  g12458(.a(n13416), .b(n13300), .O(n13546));
  invx  g12459(.a(n13546), .O(n13547));
  andx  g12460(.a(n13547), .b(n13423), .O(n13548));
  andx  g12461(.a(n13422), .b(n13298), .O(n13549));
  orx   g12462(.a(n13436), .b(n13549), .O(n13550));
  andx  g12463(.a(n13550), .b(n13548), .O(n13551));
  invx  g12464(.a(n13551), .O(n13552));
  andx  g12465(.a(n13552), .b(n13545), .O(n13553));
  andx  g12466(.a(n13543), .b(n13540), .O(n13554));
  andx  g12467(.a(n13534), .b(n13445), .O(n13555));
  orx   g12468(.a(n13555), .b(n13554), .O(n13556));
  andx  g12469(.a(n13551), .b(n13556), .O(n13557));
  orx   g12470(.a(n13557), .b(n13553), .O(po19));
  orx   g12471(.a(n13434), .b(n12962), .O(n13559));
  orx   g12472(.a(n13559), .b(n13126), .O(n13560));
  andx  g12473(.a(n13560), .b(n13288), .O(n13561));
  orx   g12474(.a(n13561), .b(n13549), .O(n13562));
  andx  g12475(.a(n13562), .b(n13548), .O(n13563));
  orx   g12476(.a(n13563), .b(n13545), .O(n13564));
  orx   g12477(.a(n13545), .b(n13549), .O(n13565));
  andx  g12478(.a(n13286), .b(n13127), .O(n13566));
  invx  g12479(.a(n13566), .O(n13567));
  orx   g12480(.a(n13567), .b(n13565), .O(n13568));
  orx   g12481(.a(n13568), .b(n12961), .O(n13569));
  andx  g12482(.a(n13569), .b(n13564), .O(n13570));
  andx  g12483(.a(n13543), .b(n13445), .O(n13571));
  invx  g12484(.a(n13571), .O(n13572));
  orx   g12485(.a(n13525), .b(n13528), .O(n13573));
  andx  g12486(.a(n13573), .b(n13452), .O(n13574));
  andx  g12487(.a(n11120), .b(n4063), .O(n13575));
  andx  g12488(.a(n13499), .b(n13501), .O(n13576));
  orx   g12489(.a(n13576), .b(n13461), .O(n13577));
  orx   g12490(.a(n13577), .b(n13575), .O(n13578));
  orx   g12491(.a(n13506), .b(n13458), .O(n13579));
  andx  g12492(.a(n13579), .b(n13502), .O(n13580));
  orx   g12493(.a(n13580), .b(n11714), .O(n13581));
  andx  g12494(.a(n13581), .b(n13578), .O(n13582));
  andx  g12495(.a(n2429), .b(n10356), .O(n13585));
  andx  g12496(.a(n2724), .b(n7902), .O(n13588));
  orx   g12497(.a(n13588), .b(n13585), .O(n13589));
  andx  g12498(.a(n11157), .b(n7902), .O(n13590));
  orx   g12499(.a(n13590), .b(n13467), .O(n13591));
  andx  g12500(.a(n13591), .b(n9470), .O(n13592));
  andx  g12501(.a(n13467), .b(n7902), .O(n13593));
  orx   g12502(.a(n13593), .b(n13592), .O(n13594));
  invx  g12503(.a(n13594), .O(n13595));
  andx  g12504(.a(n13595), .b(n13589), .O(n13596));
  invx  g12505(.a(n13596), .O(n13597));
  orx   g12506(.a(n13595), .b(n13589), .O(n13598));
  andx  g12507(.a(n13598), .b(n13597), .O(n13599));
  invx  g12508(.a(n13599), .O(n13600));
  andx  g12509(.a(n13483), .b(n13494), .O(n13601));
  invx  g12510(.a(n13601), .O(n13602));
  andx  g12511(.a(n13489), .b(n13479), .O(n13603));
  orx   g12512(.a(n13603), .b(n13490), .O(n13604));
  andx  g12513(.a(n13604), .b(n13602), .O(n13605));
  andx  g12514(.a(n10751), .b(n4114), .O(n13606));
  invx  g12515(.a(n13606), .O(n13607));
  andx  g12516(.a(n13607), .b(n13605), .O(n13608));
  orx   g12517(.a(n13483), .b(n13494), .O(n13609));
  andx  g12518(.a(n13609), .b(n13484), .O(n13610));
  orx   g12519(.a(n13610), .b(n13601), .O(n13611));
  andx  g12520(.a(n13606), .b(n13611), .O(n13612));
  orx   g12521(.a(n13612), .b(n13608), .O(n13613));
  orx   g12522(.a(n13613), .b(n13600), .O(n13614));
  orx   g12523(.a(n13606), .b(n13611), .O(n13615));
  orx   g12524(.a(n13607), .b(n13605), .O(n13616));
  andx  g12525(.a(n13616), .b(n13615), .O(n13617));
  orx   g12526(.a(n13617), .b(n13599), .O(n13618));
  andx  g12527(.a(n13618), .b(n13614), .O(n13619));
  orx   g12528(.a(n13619), .b(n13582), .O(n13620));
  invx  g12529(.a(n13575), .O(n13621));
  andx  g12530(.a(n13580), .b(n13621), .O(n13622));
  andx  g12531(.a(n13577), .b(n11120), .O(n13623));
  orx   g12532(.a(n13623), .b(n13622), .O(n13624));
  andx  g12533(.a(n13617), .b(n13599), .O(n13625));
  andx  g12534(.a(n13613), .b(n13600), .O(n13626));
  orx   g12535(.a(n13626), .b(n13625), .O(n13627));
  orx   g12536(.a(n13627), .b(n13624), .O(n13628));
  andx  g12537(.a(n13628), .b(n13620), .O(n13629));
  andx  g12538(.a(n13519), .b(n13508), .O(n13630));
  invx  g12539(.a(n13630), .O(n13631));
  orx   g12540(.a(n13506), .b(n13503), .O(n13632));
  orx   g12541(.a(n13499), .b(n13462), .O(n13633));
  andx  g12542(.a(n13633), .b(n13632), .O(n13634));
  andx  g12543(.a(n13513), .b(n13634), .O(n13635));
  orx   g12544(.a(n13635), .b(n13515), .O(n13636));
  andx  g12545(.a(n13636), .b(n13631), .O(n13637));
  andx  g12546(.a(n11451), .b(n3721), .O(n13638));
  invx  g12547(.a(n13638), .O(n13639));
  andx  g12548(.a(n13639), .b(n13637), .O(n13640));
  orx   g12549(.a(n13519), .b(n13508), .O(n13641));
  andx  g12550(.a(n13641), .b(n13514), .O(n13642));
  orx   g12551(.a(n13642), .b(n13630), .O(n13643));
  andx  g12552(.a(n13638), .b(n13643), .O(n13644));
  orx   g12553(.a(n13644), .b(n13640), .O(n13645));
  orx   g12554(.a(n13645), .b(n13629), .O(n13646));
  andx  g12555(.a(n13627), .b(n13624), .O(n13647));
  andx  g12556(.a(n13619), .b(n13582), .O(n13648));
  orx   g12557(.a(n13648), .b(n13647), .O(n13649));
  orx   g12558(.a(n13638), .b(n13643), .O(n13650));
  orx   g12559(.a(n13639), .b(n13637), .O(n13651));
  andx  g12560(.a(n13651), .b(n13650), .O(n13652));
  orx   g12561(.a(n13652), .b(n13649), .O(n13653));
  andx  g12562(.a(n13653), .b(n13646), .O(n13654));
  andx  g12563(.a(n13654), .b(n13574), .O(n13655));
  andx  g12564(.a(n13532), .b(n13449), .O(n13656));
  orx   g12565(.a(n13656), .b(n13529), .O(n13657));
  andx  g12566(.a(n13652), .b(n13649), .O(n13658));
  andx  g12567(.a(n13645), .b(n13629), .O(n13659));
  orx   g12568(.a(n13659), .b(n13658), .O(n13660));
  andx  g12569(.a(n13660), .b(n13657), .O(n13661));
  orx   g12570(.a(n13661), .b(n13655), .O(n13662));
  andx  g12571(.a(n13662), .b(n13572), .O(n13663));
  andx  g12572(.a(n13663), .b(n13570), .O(n13664));
  invx  g12573(.a(n13662), .O(n13665));
  andx  g12574(.a(n13665), .b(n13571), .O(n13666));
  andx  g12575(.a(n13426), .b(n13297), .O(n13667));
  orx   g12576(.a(n13546), .b(n13667), .O(n13668));
  andx  g12577(.a(n13286), .b(n13130), .O(n13669));
  andx  g12578(.a(n13669), .b(n13127), .O(n13670));
  orx   g12579(.a(n13670), .b(n13287), .O(n13671));
  andx  g12580(.a(n13671), .b(n13427), .O(n13672));
  orx   g12581(.a(n13672), .b(n13668), .O(n13673));
  andx  g12582(.a(n13673), .b(n13556), .O(n13674));
  andx  g12583(.a(n13556), .b(n13427), .O(n13675));
  andx  g12584(.a(n13566), .b(n13675), .O(n13676));
  andx  g12585(.a(n13676), .b(n13141), .O(n13677));
  orx   g12586(.a(n13677), .b(n13674), .O(n13678));
  andx  g12587(.a(n13665), .b(n13678), .O(n13679));
  orx   g12588(.a(n13679), .b(n13666), .O(n13680));
  orx   g12589(.a(n13680), .b(n13664), .O(po20));
  andx  g12590(.a(n13638), .b(n13649), .O(n13682));
  invx  g12591(.a(n13682), .O(n13683));
  andx  g12592(.a(n13639), .b(n13629), .O(n13684));
  orx   g12593(.a(n13684), .b(n13637), .O(n13685));
  andx  g12594(.a(n13685), .b(n13683), .O(n13686));
  andx  g12595(.a(n11451), .b(n4063), .O(n13687));
  invx  g12596(.a(n13687), .O(n13688));
  orx   g12597(.a(n13619), .b(n13622), .O(n13689));
  andx  g12598(.a(n13689), .b(n13581), .O(n13690));
  andx  g12599(.a(n13690), .b(n13688), .O(n13691));
  andx  g12600(.a(n13627), .b(n13578), .O(n13692));
  orx   g12601(.a(n13692), .b(n13623), .O(n13693));
  andx  g12602(.a(n13693), .b(n11451), .O(n13694));
  orx   g12603(.a(n13694), .b(n13691), .O(n13695));
  andx  g12604(.a(n11157), .b(n10356), .O(n13696));
  orx   g12605(.a(n13696), .b(n13594), .O(n13697));
  andx  g12606(.a(n13697), .b(n7902), .O(n13698));
  andx  g12607(.a(n13594), .b(n10356), .O(n13699));
  orx   g12608(.a(n13699), .b(n13698), .O(n13700));
  invx  g12609(.a(n13700), .O(n13701));
  andx  g12610(.a(n2724), .b(n10356), .O(n13704));
  andx  g12611(.a(n2429), .b(n10751), .O(n13707));
  orx   g12612(.a(n13707), .b(n13704), .O(n13708));
  andx  g12613(.a(n13708), .b(n13701), .O(n13709));
  invx  g12614(.a(n13709), .O(n13710));
  orx   g12615(.a(n13708), .b(n13701), .O(n13711));
  andx  g12616(.a(n13711), .b(n13710), .O(n13712));
  andx  g12617(.a(n13611), .b(n13600), .O(n13713));
  invx  g12618(.a(n13713), .O(n13714));
  andx  g12619(.a(n13605), .b(n13599), .O(n13715));
  orx   g12620(.a(n13715), .b(n13607), .O(n13716));
  andx  g12621(.a(n13716), .b(n13714), .O(n13717));
  andx  g12622(.a(n11120), .b(n4114), .O(n13718));
  invx  g12623(.a(n13718), .O(n13719));
  andx  g12624(.a(n13719), .b(n13717), .O(n13720));
  invx  g12625(.a(n13720), .O(n13721));
  orx   g12626(.a(n13719), .b(n13717), .O(n13722));
  andx  g12627(.a(n13722), .b(n13721), .O(n13723));
  andx  g12628(.a(n13723), .b(n13712), .O(n13724));
  invx  g12629(.a(n13712), .O(n13725));
  invx  g12630(.a(n13722), .O(n13726));
  orx   g12631(.a(n13726), .b(n13720), .O(n13727));
  andx  g12632(.a(n13727), .b(n13725), .O(n13728));
  orx   g12633(.a(n13728), .b(n13724), .O(n13729));
  andx  g12634(.a(n13729), .b(n13695), .O(n13730));
  orx   g12635(.a(n13693), .b(n13687), .O(n13731));
  orx   g12636(.a(n13690), .b(n12000), .O(n13732));
  andx  g12637(.a(n13732), .b(n13731), .O(n13733));
  orx   g12638(.a(n13727), .b(n13725), .O(n13734));
  orx   g12639(.a(n13723), .b(n13712), .O(n13735));
  andx  g12640(.a(n13735), .b(n13734), .O(n13736));
  andx  g12641(.a(n13736), .b(n13733), .O(n13737));
  orx   g12642(.a(n13737), .b(n13730), .O(n13738));
  andx  g12643(.a(n13738), .b(n13686), .O(n13739));
  orx   g12644(.a(n13638), .b(n13649), .O(n13740));
  andx  g12645(.a(n13740), .b(n13643), .O(n13741));
  orx   g12646(.a(n13741), .b(n13682), .O(n13742));
  orx   g12647(.a(n13736), .b(n13733), .O(n13743));
  orx   g12648(.a(n13729), .b(n13695), .O(n13744));
  andx  g12649(.a(n13744), .b(n13743), .O(n13745));
  andx  g12650(.a(n13745), .b(n13742), .O(n13746));
  orx   g12651(.a(n13746), .b(n13739), .O(n13747));
  andx  g12652(.a(n13654), .b(n13657), .O(n13748));
  orx   g12653(.a(n13748), .b(n13747), .O(n13749));
  andx  g12654(.a(n13748), .b(n13747), .O(n13750));
  invx  g12655(.a(n13750), .O(n13751));
  andx  g12656(.a(n13751), .b(n13749), .O(n13752));
  invx  g12657(.a(n13752), .O(n13753));
  andx  g12658(.a(n13572), .b(n13570), .O(n13754));
  orx   g12659(.a(n13754), .b(n13665), .O(n13755));
  orx   g12660(.a(n13755), .b(n13753), .O(n13756));
  orx   g12661(.a(n13571), .b(n13678), .O(n13757));
  andx  g12662(.a(n13757), .b(n13662), .O(n13758));
  orx   g12663(.a(n13758), .b(n13752), .O(n13759));
  andx  g12664(.a(n13759), .b(n13756), .O(po21));
  andx  g12665(.a(n13729), .b(n13731), .O(n13761));
  orx   g12666(.a(n13761), .b(n13694), .O(n13762));
  invx  g12667(.a(n13762), .O(n13763));
  andx  g12668(.a(n2429), .b(n11120), .O(n13766));
  andx  g12669(.a(n2724), .b(n10751), .O(n13769));
  orx   g12670(.a(n13769), .b(n13766), .O(n13770));
  andx  g12671(.a(n11157), .b(n10751), .O(n13771));
  orx   g12672(.a(n13771), .b(n13700), .O(n13772));
  andx  g12673(.a(n13772), .b(n10356), .O(n13773));
  andx  g12674(.a(n13700), .b(n10751), .O(n13774));
  orx   g12675(.a(n13774), .b(n13773), .O(n13775));
  invx  g12676(.a(n13775), .O(n13776));
  andx  g12677(.a(n13776), .b(n13770), .O(n13777));
  invx  g12678(.a(n13777), .O(n13778));
  orx   g12679(.a(n13776), .b(n13770), .O(n13779));
  andx  g12680(.a(n13779), .b(n13778), .O(n13780));
  invx  g12681(.a(n13780), .O(n13781));
  invx  g12682(.a(n13717), .O(n13782));
  andx  g12683(.a(n13782), .b(n13725), .O(n13783));
  invx  g12684(.a(n13783), .O(n13784));
  andx  g12685(.a(n13717), .b(n13712), .O(n13785));
  orx   g12686(.a(n13785), .b(n13719), .O(n13786));
  andx  g12687(.a(n13786), .b(n13784), .O(n13787));
  andx  g12688(.a(n11451), .b(n4114), .O(n13788));
  invx  g12689(.a(n13788), .O(n13789));
  invx  g12690(.a(n13787), .O(n13791));
  andx  g12691(.a(n13788), .b(n13791), .O(n13792));
  andx  g12692(.a(n4113), .b(n13781), .O(n13796));
  orx   g12693(.a(n13796), .b(n13788), .O(n13797));
  andx  g12694(.a(n13797), .b(n13763), .O(n13798));
  invx  g12695(.a(n13796), .O(n13799));
  andx  g12696(.a(n13799), .b(n13789), .O(n13800));
  andx  g12697(.a(n13800), .b(n13762), .O(n13801));
  orx   g12698(.a(n13801), .b(n13798), .O(n13802));
  andx  g12699(.a(n13738), .b(n13742), .O(n13803));
  andx  g12700(.a(n13803), .b(n13802), .O(n13804));
  invx  g12701(.a(n13804), .O(n13805));
  orx   g12702(.a(n13803), .b(n13802), .O(n13806));
  andx  g12703(.a(n13806), .b(n13805), .O(n13807));
  andx  g12704(.a(n13758), .b(n13749), .O(n13808));
  orx   g12705(.a(n13808), .b(n13750), .O(n13809));
  orx   g12706(.a(n13809), .b(n13807), .O(n13810));
  invx  g12707(.a(n13807), .O(n13811));
  orx   g12708(.a(n13745), .b(n13742), .O(n13812));
  orx   g12709(.a(n13738), .b(n13686), .O(n13813));
  andx  g12710(.a(n13813), .b(n13812), .O(n13814));
  orx   g12711(.a(n13660), .b(n13574), .O(n13815));
  andx  g12712(.a(n13815), .b(n13814), .O(n13816));
  andx  g12713(.a(n13756), .b(n13751), .O(n13818));
  orx   g12714(.a(n13818), .b(n13811), .O(n13819));
  andx  g12715(.a(n13819), .b(n13810), .O(po22));
  andx  g12716(.a(n13809), .b(n13806), .O(n13821));
  andx  g12717(.a(n13797), .b(n13762), .O(n13822));
  invx  g12718(.a(n13822), .O(n13823));
  andx  g12719(.a(n13823), .b(n13805), .O(n13824));
  invx  g12720(.a(n13824), .O(n13825));
  orx   g12721(.a(n13825), .b(n13821), .O(n13826));
  andx  g12722(.a(n13775), .b(n11120), .O(n13827));
  invx  g12723(.a(n13827), .O(n13828));
  andx  g12724(.a(n11157), .b(n11120), .O(n13829));
  invx  g12725(.a(n13829), .O(n13830));
  andx  g12726(.a(n13830), .b(n13776), .O(n13831));
  orx   g12727(.a(n13831), .b(n11380), .O(n13832));
  andx  g12728(.a(n13832), .b(n13828), .O(n13833));
  invx  g12729(.a(n13833), .O(n13834));
  andx  g12730(.a(n2724), .b(n11120), .O(n13837));
  andx  g12731(.a(n2429), .b(n11451), .O(n13840));
  orx   g12732(.a(n13840), .b(n13837), .O(n13841));
  andx  g12733(.a(n13841), .b(n13834), .O(n13842));
  invx  g12734(.a(n13842), .O(n13843));
  orx   g12735(.a(n13841), .b(n13834), .O(n13844));
  andx  g12736(.a(n13844), .b(n13843), .O(n13845));
  invx  g12737(.a(n13845), .O(n13846));
  andx  g12738(.a(n13788), .b(n13781), .O(n13847));
  andx  g12739(.a(n13791), .b(n13781), .O(n13848));
  orx   g12740(.a(n13848), .b(n13847), .O(n13849));
  orx   g12741(.a(n13849), .b(n13792), .O(n13850));
  andx  g12742(.a(n13850), .b(n13846), .O(n13851));
  invx  g12743(.a(n13850), .O(n13852));
  andx  g12744(.a(n13852), .b(n13845), .O(n13853));
  orx   g12745(.a(n13853), .b(n13851), .O(n13854));
  invx  g12746(.a(n13854), .O(n13855));
  andx  g12747(.a(n13855), .b(n13826), .O(n13856));
  orx   g12748(.a(n13800), .b(n13762), .O(n13857));
  orx   g12749(.a(n13797), .b(n13763), .O(n13858));
  andx  g12750(.a(n13858), .b(n13857), .O(n13859));
  invx  g12751(.a(n13803), .O(n13860));
  andx  g12752(.a(n13860), .b(n13859), .O(n13861));
  andx  g12753(.a(n13824), .b(n13819), .O(n13863));
  andx  g12754(.a(n13854), .b(n13863), .O(n13864));
  orx   g12755(.a(n13864), .b(n13856), .O(po23));
  andx  g12756(.a(n11451), .b(n2724), .O(n13866));
  invx  g12757(.a(n13866), .O(n13867));
  andx  g12758(.a(n13850), .b(n13845), .O(n13868));
  invx  g12759(.a(n13868), .O(n13869));
  andx  g12760(.a(n13869), .b(n13867), .O(n13870));
  andx  g12761(.a(n13868), .b(n13866), .O(n13871));
  orx   g12762(.a(n13871), .b(n13870), .O(n13872));
  invx  g12763(.a(n13872), .O(n13873));
  andx  g12764(.a(n13834), .b(n11120), .O(n13874));
  invx  g12765(.a(n13874), .O(n13875));
  andx  g12766(.a(n13833), .b(n13830), .O(n13876));
  orx   g12767(.a(n13876), .b(n12000), .O(n13877));
  andx  g12768(.a(n13877), .b(n13875), .O(n13878));
  invx  g12769(.a(n13878), .O(n13879));
  andx  g12770(.a(n13854), .b(n13806), .O(n13880));
  andx  g12771(.a(n13749), .b(n13662), .O(n13881));
  andx  g12772(.a(n13881), .b(n13880), .O(n13882));
  andx  g12773(.a(n13882), .b(n13678), .O(n13883));
  andx  g12774(.a(n13854), .b(n13822), .O(n13884));
  andx  g12775(.a(n13749), .b(n13571), .O(n13885));
  andx  g12776(.a(n13885), .b(n13662), .O(n13886));
  orx   g12777(.a(n13886), .b(n13750), .O(n13887));
  andx  g12778(.a(n13887), .b(n13806), .O(n13888));
  orx   g12779(.a(n13888), .b(n13804), .O(n13889));
  andx  g12780(.a(n13889), .b(n13854), .O(n13890));
  orx   g12781(.a(n13890), .b(n13884), .O(n13891));
  orx   g12782(.a(n13891), .b(n13883), .O(n13892));
  andx  g12783(.a(n13892), .b(n13879), .O(n13893));
  invx  g12784(.a(n13883), .O(n13894));
  invx  g12785(.a(n13884), .O(n13895));
  orx   g12786(.a(n13816), .b(n13572), .O(n13896));
  orx   g12787(.a(n13896), .b(n13665), .O(n13897));
  andx  g12788(.a(n13897), .b(n13751), .O(n13898));
  orx   g12789(.a(n13898), .b(n13861), .O(n13899));
  andx  g12790(.a(n13899), .b(n13805), .O(n13900));
  orx   g12791(.a(n13900), .b(n13855), .O(n13901));
  andx  g12792(.a(n13901), .b(n13895), .O(n13902));
  andx  g12793(.a(n13902), .b(n13894), .O(n13903));
  andx  g12794(.a(n13903), .b(n13878), .O(n13904));
  orx   g12795(.a(n13904), .b(n13893), .O(n13905));
  andx  g12796(.a(n13905), .b(n13873), .O(n13906));
  orx   g12797(.a(n13903), .b(n13878), .O(n13907));
  orx   g12798(.a(n13892), .b(n13879), .O(n13908));
  andx  g12799(.a(n13908), .b(n13907), .O(n13909));
  andx  g12800(.a(n13909), .b(n13872), .O(n13910));
  orx   g12801(.a(n13910), .b(n13906), .O(po24));
endmodule


