// Benchmark "top" written by ABC on Fri Feb  7 13:42:49 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22;
  wire n65, n66, n67, n68, n70, n71, n73, n74, n75, n78, n79, n81, n82, n84,
    n85, n87, n88, n90, n91, n93, n94, n96, n97, n99, n100, n102, n103,
    n105, n106, n108, n109, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n198, n199, n201, n202, n204, n205,
    n207, n208, n210, n211, n213, n214, n216, n217, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258;
  bufx g000(.A(n114), .O(n65));
  bufx g001(.A(n220), .O(n66));
  bufx g002(.A(n220), .O(n67));
  bufx g003(.A(n220), .O(n68));
  bufx g004(.A(n220), .O(po22));
  bufx g005(.A(n112), .O(n70));
  invx g006(.A(n222), .O(n71));
  invx g007(.A(n71), .O(po21));
  invx g008(.A(n71), .O(n73));
  invx g009(.A(n71), .O(n74));
  invx g010(.A(n71), .O(n75));
  xorx g011(.A(pi41), .B(pi40), .O(po20));
  orx  g012(.A(n79), .B(n78), .O(po19));
  andx g013(.A(pi39), .B(n66), .O(n78));
  andx g014(.A(pi38), .B(n73), .O(n79));
  orx  g015(.A(n82), .B(n81), .O(po18));
  andx g016(.A(pi37), .B(n67), .O(n81));
  andx g017(.A(pi36), .B(n74), .O(n82));
  orx  g018(.A(n85), .B(n84), .O(po17));
  andx g019(.A(pi35), .B(n68), .O(n84));
  andx g020(.A(pi34), .B(n75), .O(n85));
  orx  g021(.A(n88), .B(n87), .O(po16));
  andx g022(.A(pi33), .B(po22), .O(n87));
  andx g023(.A(pi32), .B(po21), .O(n88));
  orx  g024(.A(n91), .B(n90), .O(po15));
  andx g025(.A(n70), .B(n189), .O(n90));
  andx g026(.A(n193), .B(n65), .O(n91));
  orx  g027(.A(n94), .B(n93), .O(po14));
  andx g028(.A(n70), .B(n120), .O(n93));
  andx g029(.A(n185), .B(n65), .O(n94));
  orx  g030(.A(n97), .B(n96), .O(po13));
  andx g031(.A(n70), .B(n177), .O(n96));
  andx g032(.A(n181), .B(n65), .O(n97));
  orx  g033(.A(n100), .B(n99), .O(po12));
  andx g034(.A(n70), .B(n169), .O(n99));
  andx g035(.A(n173), .B(n65), .O(n100));
  orx  g036(.A(n103), .B(n102), .O(po11));
  andx g037(.A(n112), .B(n161), .O(n102));
  andx g038(.A(n165), .B(n65), .O(n103));
  orx  g039(.A(n106), .B(n105), .O(po10));
  andx g040(.A(n112), .B(n153), .O(n105));
  andx g041(.A(n157), .B(n65), .O(n106));
  orx  g042(.A(n109), .B(n108), .O(po09));
  andx g043(.A(n112), .B(n142), .O(n108));
  andx g044(.A(n146), .B(n114), .O(n109));
  orx  g045(.A(n113), .B(n111), .O(po08));
  andx g046(.A(n112), .B(n149), .O(n111));
  invx g047(.A(n114), .O(n112));
  andx g048(.A(n194), .B(n114), .O(n113));
  orx  g049(.A(n116), .B(n115), .O(n114));
  andx g050(.A(n192), .B(n189), .O(n115));
  andx g051(.A(n118), .B(n117), .O(n116));
  orx  g052(.A(n184), .B(n124), .O(n117));
  andx g053(.A(n188), .B(n119), .O(n118));
  orx  g054(.A(n123), .B(n120), .O(n119));
  orx  g055(.A(n122), .B(n121), .O(n120));
  andx g056(.A(pi31), .B(n66), .O(n121));
  andx g057(.A(pi24), .B(n73), .O(n122));
  andx g058(.A(n184), .B(n124), .O(n123));
  orx  g059(.A(n126), .B(n125), .O(n124));
  andx g060(.A(n180), .B(n177), .O(n125));
  andx g061(.A(n176), .B(n127), .O(n126));
  orx  g062(.A(n129), .B(n128), .O(n127));
  andx g063(.A(n172), .B(n169), .O(n128));
  andx g064(.A(n168), .B(n130), .O(n129));
  orx  g065(.A(n132), .B(n131), .O(n130));
  andx g066(.A(n164), .B(n161), .O(n131));
  andx g067(.A(n160), .B(n133), .O(n132));
  orx  g068(.A(n135), .B(n134), .O(n133));
  andx g069(.A(n156), .B(n153), .O(n134));
  andx g070(.A(n152), .B(n136), .O(n135));
  orx  g071(.A(n138), .B(n137), .O(n136));
  andx g072(.A(n145), .B(n142), .O(n137));
  andx g073(.A(n140), .B(n139), .O(n138));
  invx g074(.A(n194), .O(n139));
  andx g075(.A(n149), .B(n141), .O(n140));
  orx  g076(.A(n145), .B(n142), .O(n141));
  orx  g077(.A(n144), .B(n143), .O(n142));
  andx g078(.A(pi07), .B(n67), .O(n143));
  andx g079(.A(pi04), .B(n74), .O(n144));
  invx g080(.A(n146), .O(n145));
  orx  g081(.A(n148), .B(n147), .O(n146));
  andx g082(.A(pi06), .B(n68), .O(n147));
  andx g083(.A(pi05), .B(n75), .O(n148));
  orx  g084(.A(n151), .B(n150), .O(n149));
  andx g085(.A(pi01), .B(po22), .O(n150));
  andx g086(.A(pi00), .B(po21), .O(n151));
  orx  g087(.A(n156), .B(n153), .O(n152));
  orx  g088(.A(n155), .B(n154), .O(n153));
  andx g089(.A(pi11), .B(n66), .O(n154));
  andx g090(.A(pi08), .B(n73), .O(n155));
  invx g091(.A(n157), .O(n156));
  orx  g092(.A(n159), .B(n158), .O(n157));
  andx g093(.A(pi10), .B(n67), .O(n158));
  andx g094(.A(pi09), .B(n74), .O(n159));
  orx  g095(.A(n164), .B(n161), .O(n160));
  orx  g096(.A(n163), .B(n162), .O(n161));
  andx g097(.A(pi15), .B(n68), .O(n162));
  andx g098(.A(pi12), .B(n75), .O(n163));
  invx g099(.A(n165), .O(n164));
  orx  g100(.A(n167), .B(n166), .O(n165));
  andx g101(.A(pi14), .B(po22), .O(n166));
  andx g102(.A(pi13), .B(po21), .O(n167));
  orx  g103(.A(n172), .B(n169), .O(n168));
  orx  g104(.A(n171), .B(n170), .O(n169));
  andx g105(.A(pi19), .B(n66), .O(n170));
  andx g106(.A(pi16), .B(n73), .O(n171));
  invx g107(.A(n173), .O(n172));
  orx  g108(.A(n175), .B(n174), .O(n173));
  andx g109(.A(pi18), .B(n67), .O(n174));
  andx g110(.A(pi17), .B(n74), .O(n175));
  orx  g111(.A(n180), .B(n177), .O(n176));
  orx  g112(.A(n179), .B(n178), .O(n177));
  andx g113(.A(pi23), .B(n68), .O(n178));
  andx g114(.A(pi20), .B(n75), .O(n179));
  invx g115(.A(n181), .O(n180));
  orx  g116(.A(n183), .B(n182), .O(n181));
  andx g117(.A(pi22), .B(po22), .O(n182));
  andx g118(.A(pi21), .B(po21), .O(n183));
  invx g119(.A(n185), .O(n184));
  orx  g120(.A(n187), .B(n186), .O(n185));
  andx g121(.A(pi28), .B(n66), .O(n186));
  andx g122(.A(pi26), .B(n73), .O(n187));
  orx  g123(.A(n192), .B(n189), .O(n188));
  orx  g124(.A(n191), .B(n190), .O(n189));
  andx g125(.A(pi30), .B(n67), .O(n190));
  andx g126(.A(pi25), .B(n74), .O(n191));
  invx g127(.A(n193), .O(n192));
  orx  g128(.A(pi29), .B(pi27), .O(n193));
  orx  g129(.A(n196), .B(n195), .O(n194));
  andx g130(.A(pi03), .B(n68), .O(n195));
  andx g131(.A(pi02), .B(n75), .O(n196));
  orx  g132(.A(n199), .B(n198), .O(po07));
  andx g133(.A(pi27), .B(po22), .O(n198));
  andx g134(.A(pi29), .B(po21), .O(n199));
  orx  g135(.A(n202), .B(n201), .O(po06));
  andx g136(.A(pi26), .B(n66), .O(n201));
  andx g137(.A(pi28), .B(n73), .O(n202));
  orx  g138(.A(n205), .B(n204), .O(po05));
  andx g139(.A(pi21), .B(n67), .O(n204));
  andx g140(.A(pi22), .B(n74), .O(n205));
  orx  g141(.A(n208), .B(n207), .O(po04));
  andx g142(.A(pi17), .B(n68), .O(n207));
  andx g143(.A(pi18), .B(n75), .O(n208));
  orx  g144(.A(n211), .B(n210), .O(po03));
  andx g145(.A(pi13), .B(po22), .O(n210));
  andx g146(.A(pi14), .B(po21), .O(n211));
  orx  g147(.A(n214), .B(n213), .O(po02));
  andx g148(.A(pi09), .B(n66), .O(n213));
  andx g149(.A(pi10), .B(n73), .O(n214));
  orx  g150(.A(n217), .B(n216), .O(po01));
  andx g151(.A(pi05), .B(n67), .O(n216));
  andx g152(.A(pi06), .B(n74), .O(n217));
  orx  g153(.A(n221), .B(n219), .O(po00));
  andx g154(.A(pi02), .B(n68), .O(n219));
  invx g155(.A(po21), .O(n220));
  andx g156(.A(pi03), .B(n75), .O(n221));
  orx  g157(.A(n224), .B(n223), .O(n222));
  andx g158(.A(pi27), .B(n258), .O(n223));
  andx g159(.A(n226), .B(n225), .O(n224));
  orx  g160(.A(n230), .B(n229), .O(n225));
  andx g161(.A(n257), .B(n227), .O(n226));
  orx  g162(.A(n228), .B(pi26), .O(n227));
  andx g163(.A(n230), .B(n229), .O(n228));
  invx g164(.A(pi28), .O(n229));
  orx  g165(.A(n232), .B(n231), .O(n230));
  andx g166(.A(n235), .B(n234), .O(n231));
  andx g167(.A(pi21), .B(n233), .O(n232));
  orx  g168(.A(n235), .B(n234), .O(n233));
  invx g169(.A(pi22), .O(n234));
  orx  g170(.A(n237), .B(n236), .O(n235));
  andx g171(.A(n240), .B(n239), .O(n236));
  andx g172(.A(pi17), .B(n238), .O(n237));
  orx  g173(.A(n240), .B(n239), .O(n238));
  invx g174(.A(pi18), .O(n239));
  orx  g175(.A(n242), .B(n241), .O(n240));
  andx g176(.A(n245), .B(n244), .O(n241));
  andx g177(.A(pi13), .B(n243), .O(n242));
  orx  g178(.A(n245), .B(n244), .O(n243));
  invx g179(.A(pi14), .O(n244));
  orx  g180(.A(n247), .B(n246), .O(n245));
  andx g181(.A(n250), .B(n249), .O(n246));
  andx g182(.A(pi09), .B(n248), .O(n247));
  orx  g183(.A(n250), .B(n249), .O(n248));
  invx g184(.A(pi10), .O(n249));
  orx  g185(.A(n252), .B(n251), .O(n250));
  andx g186(.A(pi05), .B(n256), .O(n251));
  andx g187(.A(n253), .B(pi02), .O(n252));
  andx g188(.A(n255), .B(n254), .O(n253));
  invx g189(.A(pi03), .O(n254));
  orx  g190(.A(pi05), .B(n256), .O(n255));
  invx g191(.A(pi06), .O(n256));
  orx  g192(.A(pi27), .B(n258), .O(n257));
  invx g193(.A(pi29), .O(n258));
endmodule


