// Benchmark "top" written by ABC on Fri Feb  7 13:47:33 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
    n48, n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n62, n63, n64,
    n65, n66, n67, n69, n70, n71, n72, n73, n74, n76, n77, n78, n79, n80,
    n81, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n364, n365, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702;
  bufx g000(.A(n507), .O(po04));
  bufx g001(.A(n582), .O(n33));
  bufx g002(.A(n272), .O(n34));
  bufx g003(.A(n436), .O(po02));
  bufx g004(.A(n556), .O(n36));
  bufx g005(.A(n453), .O(n37));
  bufx g006(.A(n100), .O(n38));
  bufx g007(.A(n192), .O(n39));
  bufx g008(.A(n683), .O(n40));
  bufx g009(.A(n683), .O(n41));
  bufx g010(.A(n540), .O(n42));
  bufx g011(.A(n101), .O(n43));
  invx g012(.A(pi01), .O(n44));
  invx g013(.A(pi01), .O(n45));
  bufx g014(.A(n702), .O(n46));
  bufx g015(.A(n702), .O(n47));
  bufx g016(.A(n702), .O(n48));
  orx  g017(.A(n51), .B(n50), .O(po15));
  andx g018(.A(n38), .B(n188), .O(n50));
  andx g019(.A(n52), .B(n43), .O(n51));
  andx g020(.A(n53), .B(n104), .O(n52));
  invx g021(.A(n184), .O(n53));
  orx  g022(.A(n56), .B(n55), .O(po13));
  andx g023(.A(n38), .B(n177), .O(n55));
  andx g024(.A(n57), .B(n43), .O(n56));
  orx  g025(.A(n59), .B(n58), .O(n57));
  andx g026(.A(n173), .B(n106), .O(n58));
  invx g027(.A(n60), .O(n59));
  orx  g028(.A(n106), .B(n173), .O(n60));
  orx  g029(.A(n63), .B(n62), .O(po11));
  andx g030(.A(n100), .B(n165), .O(n62));
  andx g031(.A(n64), .B(n43), .O(n63));
  orx  g032(.A(n66), .B(n65), .O(n64));
  andx g033(.A(n161), .B(n108), .O(n65));
  invx g034(.A(n67), .O(n66));
  orx  g035(.A(n108), .B(n161), .O(n67));
  orx  g036(.A(n70), .B(n69), .O(po09));
  andx g037(.A(n100), .B(n153), .O(n69));
  andx g038(.A(n71), .B(n43), .O(n70));
  orx  g039(.A(n73), .B(n72), .O(n71));
  andx g040(.A(n149), .B(n110), .O(n72));
  invx g041(.A(n74), .O(n73));
  orx  g042(.A(n110), .B(n149), .O(n74));
  orx  g043(.A(n77), .B(n76), .O(po07));
  andx g044(.A(n100), .B(n141), .O(n76));
  andx g045(.A(n78), .B(n43), .O(n77));
  orx  g046(.A(n80), .B(n79), .O(n78));
  andx g047(.A(n137), .B(n112), .O(n79));
  invx g048(.A(n81), .O(n80));
  orx  g049(.A(n112), .B(n137), .O(n81));
  orx  g050(.A(n84), .B(n83), .O(po05));
  andx g051(.A(n100), .B(n130), .O(n83));
  andx g052(.A(n85), .B(n43), .O(n84));
  orx  g053(.A(n87), .B(n86), .O(n85));
  andx g054(.A(n126), .B(n114), .O(n86));
  invx g055(.A(n88), .O(n87));
  orx  g056(.A(n114), .B(n126), .O(n88));
  orx  g057(.A(n94), .B(n90), .O(po03));
  andx g058(.A(n91), .B(n43), .O(n90));
  andx g059(.A(n93), .B(n92), .O(n91));
  orx  g060(.A(n398), .B(n117), .O(n92));
  invx g061(.A(n116), .O(n93));
  andx g062(.A(n100), .B(n121), .O(n94));
  orx  g063(.A(n98), .B(n96), .O(po01));
  invx g064(.A(n97), .O(n96));
  orx  g065(.A(n38), .B(n398), .O(n97));
  andx g066(.A(pi00), .B(n99), .O(n98));
  orx  g067(.A(n100), .B(n44), .O(n99));
  invx g068(.A(n101), .O(n100));
  orx  g069(.A(n103), .B(n102), .O(n101));
  andx g070(.A(n188), .B(n694), .O(n102));
  andx g071(.A(n184), .B(n104), .O(n103));
  orx  g072(.A(n105), .B(n174), .O(n104));
  andx g073(.A(n172), .B(n106), .O(n105));
  orx  g074(.A(n107), .B(n162), .O(n106));
  andx g075(.A(n160), .B(n108), .O(n107));
  orx  g076(.A(n109), .B(n150), .O(n108));
  andx g077(.A(n148), .B(n110), .O(n109));
  orx  g078(.A(n111), .B(n138), .O(n110));
  andx g079(.A(n136), .B(n112), .O(n111));
  orx  g080(.A(n113), .B(n127), .O(n112));
  andx g081(.A(n125), .B(n114), .O(n113));
  orx  g082(.A(n116), .B(n115), .O(n114));
  andx g083(.A(n121), .B(n46), .O(n115));
  andx g084(.A(n398), .B(n117), .O(n116));
  orx  g085(.A(n120), .B(n118), .O(n117));
  andx g086(.A(n119), .B(n48), .O(n118));
  invx g087(.A(n121), .O(n119));
  andx g088(.A(pi03), .B(n121), .O(n120));
  orx  g089(.A(n123), .B(n122), .O(n121));
  andx g090(.A(n404), .B(n39), .O(n122));
  andx g091(.A(pi02), .B(n124), .O(n123));
  orx  g092(.A(n190), .B(n45), .O(n124));
  invx g093(.A(n126), .O(n125));
  orx  g094(.A(n128), .B(n127), .O(n126));
  andx g095(.A(n130), .B(n40), .O(n127));
  andx g096(.A(n129), .B(pi05), .O(n128));
  invx g097(.A(n130), .O(n129));
  orx  g098(.A(n135), .B(n131), .O(n130));
  andx g099(.A(n132), .B(n39), .O(n131));
  andx g100(.A(n134), .B(n133), .O(n132));
  orx  g101(.A(n37), .B(n208), .O(n133));
  orx  g102(.A(n404), .B(n209), .O(n134));
  andx g103(.A(n190), .B(n213), .O(n135));
  invx g104(.A(n137), .O(n136));
  orx  g105(.A(n139), .B(n138), .O(n137));
  andx g106(.A(n141), .B(n42), .O(n138));
  andx g107(.A(n140), .B(pi07), .O(n139));
  invx g108(.A(n141), .O(n140));
  orx  g109(.A(n143), .B(n142), .O(n141));
  andx g110(.A(n190), .B(n222), .O(n142));
  andx g111(.A(n144), .B(n39), .O(n143));
  orx  g112(.A(n146), .B(n145), .O(n144));
  andx g113(.A(n218), .B(n205), .O(n145));
  invx g114(.A(n147), .O(n146));
  orx  g115(.A(n205), .B(n218), .O(n147));
  invx g116(.A(n149), .O(n148));
  orx  g117(.A(n151), .B(n150), .O(n149));
  andx g118(.A(n153), .B(n523), .O(n150));
  andx g119(.A(n152), .B(pi09), .O(n151));
  invx g120(.A(n153), .O(n152));
  orx  g121(.A(n155), .B(n154), .O(n153));
  andx g122(.A(n190), .B(n233), .O(n154));
  andx g123(.A(n156), .B(n39), .O(n155));
  orx  g124(.A(n158), .B(n157), .O(n156));
  andx g125(.A(n229), .B(n203), .O(n157));
  invx g126(.A(n159), .O(n158));
  orx  g127(.A(n203), .B(n229), .O(n159));
  invx g128(.A(n161), .O(n160));
  orx  g129(.A(n163), .B(n162), .O(n161));
  andx g130(.A(n165), .B(n695), .O(n162));
  andx g131(.A(n164), .B(pi11), .O(n163));
  invx g132(.A(n165), .O(n164));
  orx  g133(.A(n167), .B(n166), .O(n165));
  andx g134(.A(n190), .B(n245), .O(n166));
  andx g135(.A(n168), .B(n39), .O(n167));
  orx  g136(.A(n170), .B(n169), .O(n168));
  andx g137(.A(n241), .B(n201), .O(n169));
  invx g138(.A(n171), .O(n170));
  orx  g139(.A(n201), .B(n241), .O(n171));
  invx g140(.A(n173), .O(n172));
  orx  g141(.A(n175), .B(n174), .O(n173));
  andx g142(.A(n177), .B(n693), .O(n174));
  andx g143(.A(n176), .B(pi13), .O(n175));
  invx g144(.A(n177), .O(n176));
  orx  g145(.A(n179), .B(n178), .O(n177));
  andx g146(.A(n190), .B(n256), .O(n178));
  andx g147(.A(n180), .B(n192), .O(n179));
  orx  g148(.A(n182), .B(n181), .O(n180));
  andx g149(.A(n252), .B(n199), .O(n181));
  invx g150(.A(n183), .O(n182));
  orx  g151(.A(n199), .B(n252), .O(n183));
  andx g152(.A(n187), .B(n185), .O(n184));
  orx  g153(.A(n186), .B(pi15), .O(n185));
  invx g154(.A(n188), .O(n186));
  orx  g155(.A(n694), .B(n188), .O(n187));
  orx  g156(.A(n191), .B(n189), .O(n188));
  andx g157(.A(n190), .B(n268), .O(n189));
  invx g158(.A(n192), .O(n190));
  andx g159(.A(n196), .B(n192), .O(n191));
  orx  g160(.A(n194), .B(n193), .O(n192));
  andx g161(.A(n692), .B(n268), .O(n193));
  andx g162(.A(n195), .B(n264), .O(n194));
  andx g163(.A(n197), .B(n694), .O(n195));
  andx g164(.A(n263), .B(n197), .O(n196));
  orx  g165(.A(n198), .B(n253), .O(n197));
  andx g166(.A(n251), .B(n199), .O(n198));
  orx  g167(.A(n200), .B(n242), .O(n199));
  andx g168(.A(n240), .B(n201), .O(n200));
  orx  g169(.A(n202), .B(n230), .O(n201));
  andx g170(.A(n228), .B(n203), .O(n202));
  orx  g171(.A(n204), .B(n219), .O(n203));
  andx g172(.A(n217), .B(n205), .O(n204));
  orx  g173(.A(n207), .B(n206), .O(n205));
  andx g174(.A(n213), .B(n47), .O(n206));
  andx g175(.A(n208), .B(n37), .O(n207));
  invx g176(.A(n209), .O(n208));
  andx g177(.A(n211), .B(n210), .O(n209));
  orx  g178(.A(n213), .B(pi03), .O(n210));
  orx  g179(.A(n48), .B(n212), .O(n211));
  invx g180(.A(n213), .O(n212));
  orx  g181(.A(n215), .B(n214), .O(n213));
  andx g182(.A(n473), .B(n34), .O(n214));
  andx g183(.A(pi04), .B(n216), .O(n215));
  orx  g184(.A(n270), .B(n45), .O(n216));
  invx g185(.A(n218), .O(n217));
  orx  g186(.A(n220), .B(n219), .O(n218));
  andx g187(.A(n222), .B(n41), .O(n219));
  andx g188(.A(n221), .B(pi05), .O(n220));
  invx g189(.A(n222), .O(n221));
  orx  g190(.A(n227), .B(n223), .O(n222));
  andx g191(.A(n224), .B(n34), .O(n223));
  andx g192(.A(n226), .B(n225), .O(n224));
  orx  g193(.A(n36), .B(n301), .O(n225));
  orx  g194(.A(n473), .B(n302), .O(n226));
  andx g195(.A(n270), .B(n306), .O(n227));
  invx g196(.A(n229), .O(n228));
  orx  g197(.A(n231), .B(n230), .O(n229));
  andx g198(.A(n233), .B(n42), .O(n230));
  andx g199(.A(n232), .B(pi07), .O(n231));
  invx g200(.A(n233), .O(n232));
  orx  g201(.A(n235), .B(n234), .O(n233));
  andx g202(.A(n270), .B(n315), .O(n234));
  andx g203(.A(n236), .B(n34), .O(n235));
  orx  g204(.A(n238), .B(n237), .O(n236));
  andx g205(.A(n311), .B(n298), .O(n237));
  invx g206(.A(n239), .O(n238));
  orx  g207(.A(n298), .B(n311), .O(n239));
  invx g208(.A(n241), .O(n240));
  orx  g209(.A(n243), .B(n242), .O(n241));
  andx g210(.A(n245), .B(n523), .O(n242));
  andx g211(.A(n244), .B(pi09), .O(n243));
  invx g212(.A(n245), .O(n244));
  orx  g213(.A(n250), .B(n246), .O(n245));
  andx g214(.A(n247), .B(n34), .O(n246));
  andx g215(.A(n249), .B(n248), .O(n247));
  orx  g216(.A(n283), .B(n296), .O(n248));
  invx g217(.A(n282), .O(n249));
  andx g218(.A(n270), .B(n287), .O(n250));
  invx g219(.A(n252), .O(n251));
  orx  g220(.A(n254), .B(n253), .O(n252));
  andx g221(.A(n256), .B(n695), .O(n253));
  andx g222(.A(n255), .B(pi11), .O(n254));
  invx g223(.A(n256), .O(n255));
  orx  g224(.A(n258), .B(n257), .O(n256));
  andx g225(.A(n270), .B(n325), .O(n257));
  andx g226(.A(n259), .B(n34), .O(n258));
  orx  g227(.A(n261), .B(n260), .O(n259));
  andx g228(.A(n321), .B(n280), .O(n260));
  invx g229(.A(n262), .O(n261));
  orx  g230(.A(n280), .B(n321), .O(n262));
  invx g231(.A(n264), .O(n263));
  andx g232(.A(n267), .B(n265), .O(n264));
  orx  g233(.A(n266), .B(pi13), .O(n265));
  invx g234(.A(n268), .O(n266));
  orx  g235(.A(n268), .B(n693), .O(n267));
  orx  g236(.A(n271), .B(n269), .O(n268));
  andx g237(.A(n270), .B(n337), .O(n269));
  invx g238(.A(n34), .O(n270));
  andx g239(.A(n277), .B(n34), .O(n271));
  orx  g240(.A(n274), .B(n273), .O(n272));
  andx g241(.A(n691), .B(n337), .O(n273));
  andx g242(.A(n276), .B(n275), .O(n274));
  invx g243(.A(n335), .O(n275));
  andx g244(.A(n692), .B(n278), .O(n276));
  andx g245(.A(n335), .B(n278), .O(n277));
  orx  g246(.A(n279), .B(n322), .O(n278));
  andx g247(.A(n320), .B(n280), .O(n279));
  orx  g248(.A(n282), .B(n281), .O(n280));
  andx g249(.A(n287), .B(n42), .O(n281));
  andx g250(.A(n296), .B(n283), .O(n282));
  orx  g251(.A(n286), .B(n284), .O(n283));
  andx g252(.A(n285), .B(n42), .O(n284));
  invx g253(.A(n287), .O(n285));
  andx g254(.A(pi07), .B(n287), .O(n286));
  orx  g255(.A(n291), .B(n288), .O(n287));
  andx g256(.A(n600), .B(n289), .O(n288));
  orx  g257(.A(n290), .B(n342), .O(n289));
  andx g258(.A(n293), .B(n40), .O(n290));
  andx g259(.A(n292), .B(n341), .O(n291));
  andx g260(.A(n293), .B(n589), .O(n292));
  orx  g261(.A(n294), .B(n591), .O(n293));
  andx g262(.A(n295), .B(n597), .O(n294));
  invx g263(.A(n359), .O(n295));
  orx  g264(.A(n297), .B(n312), .O(n296));
  andx g265(.A(n310), .B(n298), .O(n297));
  orx  g266(.A(n300), .B(n299), .O(n298));
  andx g267(.A(n306), .B(n46), .O(n299));
  andx g268(.A(n301), .B(n36), .O(n300));
  invx g269(.A(n302), .O(n301));
  andx g270(.A(n304), .B(n303), .O(n302));
  orx  g271(.A(n306), .B(pi03), .O(n303));
  orx  g272(.A(n47), .B(n305), .O(n304));
  invx g273(.A(n306), .O(n305));
  orx  g274(.A(n308), .B(n307), .O(n306));
  andx g275(.A(n341), .B(n577), .O(n307));
  andx g276(.A(pi06), .B(n309), .O(n308));
  orx  g277(.A(n701), .B(n342), .O(n309));
  invx g278(.A(n311), .O(n310));
  orx  g279(.A(n313), .B(n312), .O(n311));
  andx g280(.A(n315), .B(n41), .O(n312));
  andx g281(.A(n314), .B(pi05), .O(n313));
  invx g282(.A(n315), .O(n314));
  orx  g283(.A(n318), .B(n316), .O(n315));
  andx g284(.A(n317), .B(n573), .O(n316));
  andx g285(.A(n341), .B(n575), .O(n317));
  andx g286(.A(n319), .B(n593), .O(n318));
  orx  g287(.A(n342), .B(n696), .O(n319));
  invx g288(.A(n321), .O(n320));
  orx  g289(.A(n323), .B(n322), .O(n321));
  andx g290(.A(n325), .B(n523), .O(n322));
  andx g291(.A(n324), .B(pi09), .O(n323));
  invx g292(.A(n325), .O(n324));
  orx  g293(.A(n334), .B(n326), .O(n325));
  andx g294(.A(n327), .B(n341), .O(n326));
  andx g295(.A(n330), .B(n328), .O(n327));
  invx g296(.A(n329), .O(n328));
  andx g297(.A(n358), .B(n331), .O(n329));
  orx  g298(.A(n331), .B(n358), .O(n330));
  andx g299(.A(n351), .B(n332), .O(n331));
  orx  g300(.A(pi07), .B(n333), .O(n332));
  invx g301(.A(n352), .O(n333));
  andx g302(.A(n352), .B(n342), .O(n334));
  andx g303(.A(n338), .B(n336), .O(n335));
  orx  g304(.A(n337), .B(pi11), .O(n336));
  invx g305(.A(n339), .O(n337));
  orx  g306(.A(n695), .B(n339), .O(n338));
  andx g307(.A(n346), .B(n340), .O(n339));
  orx  g308(.A(n361), .B(n341), .O(n340));
  invx g309(.A(n342), .O(n341));
  orx  g310(.A(n343), .B(n690), .O(n342));
  andx g311(.A(n360), .B(n344), .O(n343));
  orx  g312(.A(n347), .B(n345), .O(n344));
  andx g313(.A(pi09), .B(n361), .O(n345));
  orx  g314(.A(n360), .B(n347), .O(n346));
  invx g315(.A(n348), .O(n347));
  orx  g316(.A(n350), .B(n349), .O(n348));
  andx g317(.A(n352), .B(n540), .O(n349));
  andx g318(.A(n358), .B(n351), .O(n350));
  orx  g319(.A(n540), .B(n352), .O(n351));
  orx  g320(.A(n356), .B(n353), .O(n352));
  andx g321(.A(n634), .B(n354), .O(n353));
  orx  g322(.A(n355), .B(n625), .O(n354));
  andx g323(.A(n618), .B(n40), .O(n355));
  andx g324(.A(n357), .B(po08), .O(n356));
  andx g325(.A(n618), .B(n631), .O(n357));
  orx  g326(.A(n359), .B(n590), .O(n358));
  andx g327(.A(n40), .B(n600), .O(n359));
  orx  g328(.A(pi09), .B(n361), .O(n360));
  andx g329(.A(n362), .B(n623), .O(n361));
  orx  g330(.A(n653), .B(n628), .O(n362));
  andx g331(.A(n364), .B(n682), .O(po14));
  andx g332(.A(n685), .B(n365), .O(n364));
  orx  g333(.A(pi14), .B(n44), .O(n365));
  orx  g334(.A(n368), .B(n367), .O(po00));
  andx g335(.A(n434), .B(n370), .O(n367));
  andx g336(.A(n369), .B(n694), .O(n368));
  orx  g337(.A(n434), .B(n370), .O(n369));
  orx  g338(.A(n372), .B(n371), .O(n370));
  andx g339(.A(n427), .B(n374), .O(n371));
  andx g340(.A(n373), .B(n693), .O(n372));
  orx  g341(.A(n427), .B(n374), .O(n373));
  orx  g342(.A(n376), .B(n375), .O(n374));
  andx g343(.A(n420), .B(n378), .O(n375));
  andx g344(.A(n377), .B(n695), .O(n376));
  orx  g345(.A(n420), .B(n378), .O(n377));
  orx  g346(.A(n380), .B(n379), .O(n378));
  andx g347(.A(n413), .B(n382), .O(n379));
  andx g348(.A(n381), .B(n523), .O(n380));
  orx  g349(.A(n413), .B(n382), .O(n381));
  orx  g350(.A(n384), .B(n383), .O(n382));
  andx g351(.A(n406), .B(n386), .O(n383));
  andx g352(.A(n385), .B(n540), .O(n384));
  orx  g353(.A(n406), .B(n386), .O(n385));
  orx  g354(.A(n388), .B(n387), .O(n386));
  andx g355(.A(n399), .B(n390), .O(n387));
  andx g356(.A(n389), .B(n41), .O(n388));
  orx  g357(.A(n399), .B(n390), .O(n389));
  orx  g358(.A(n392), .B(n391), .O(n390));
  andx g359(.A(n394), .B(n398), .O(n391));
  andx g360(.A(n393), .B(n48), .O(n392));
  orx  g361(.A(n398), .B(n394), .O(n393));
  orx  g362(.A(n396), .B(n395), .O(n394));
  andx g363(.A(n404), .B(po02), .O(n395));
  andx g364(.A(pi02), .B(n397), .O(n396));
  orx  g365(.A(n435), .B(n45), .O(n397));
  orx  g366(.A(pi00), .B(n701), .O(n398));
  orx  g367(.A(n405), .B(n400), .O(n399));
  andx g368(.A(n401), .B(po02), .O(n400));
  andx g369(.A(n403), .B(n402), .O(n401));
  orx  g370(.A(n37), .B(n454), .O(n402));
  orx  g371(.A(n404), .B(n455), .O(n403));
  invx g372(.A(n37), .O(n404));
  andx g373(.A(n459), .B(n435), .O(n405));
  orx  g374(.A(n408), .B(n407), .O(n406));
  andx g375(.A(n468), .B(n435), .O(n407));
  andx g376(.A(n409), .B(po02), .O(n408));
  orx  g377(.A(n411), .B(n410), .O(n409));
  andx g378(.A(n464), .B(n450), .O(n410));
  invx g379(.A(n412), .O(n411));
  orx  g380(.A(n450), .B(n464), .O(n412));
  orx  g381(.A(n415), .B(n414), .O(n413));
  andx g382(.A(n480), .B(n435), .O(n414));
  andx g383(.A(n416), .B(po02), .O(n415));
  orx  g384(.A(n418), .B(n417), .O(n416));
  andx g385(.A(n476), .B(n448), .O(n417));
  invx g386(.A(n419), .O(n418));
  orx  g387(.A(n448), .B(n476), .O(n419));
  orx  g388(.A(n422), .B(n421), .O(n420));
  andx g389(.A(n492), .B(n435), .O(n421));
  andx g390(.A(n423), .B(po02), .O(n422));
  orx  g391(.A(n425), .B(n424), .O(n423));
  andx g392(.A(n488), .B(n446), .O(n424));
  invx g393(.A(n426), .O(n425));
  orx  g394(.A(n446), .B(n488), .O(n426));
  orx  g395(.A(n429), .B(n428), .O(n427));
  andx g396(.A(n503), .B(n435), .O(n428));
  andx g397(.A(n430), .B(po02), .O(n429));
  orx  g398(.A(n432), .B(n431), .O(n430));
  andx g399(.A(n499), .B(n444), .O(n431));
  invx g400(.A(n433), .O(n432));
  orx  g401(.A(n444), .B(n499), .O(n433));
  andx g402(.A(n435), .B(n440), .O(n434));
  invx g403(.A(po02), .O(n435));
  orx  g404(.A(n438), .B(n437), .O(n436));
  andx g405(.A(n692), .B(n440), .O(n437));
  andx g406(.A(n441), .B(n439), .O(n438));
  orx  g407(.A(n440), .B(n693), .O(n439));
  andx g408(.A(n505), .B(n515), .O(n440));
  andx g409(.A(n442), .B(n694), .O(n441));
  orx  g410(.A(n443), .B(n500), .O(n442));
  andx g411(.A(n498), .B(n444), .O(n443));
  orx  g412(.A(n445), .B(n489), .O(n444));
  andx g413(.A(n487), .B(n446), .O(n445));
  orx  g414(.A(n447), .B(n477), .O(n446));
  andx g415(.A(n475), .B(n448), .O(n447));
  orx  g416(.A(n449), .B(n465), .O(n448));
  andx g417(.A(n463), .B(n450), .O(n449));
  orx  g418(.A(n452), .B(n451), .O(n450));
  andx g419(.A(n459), .B(n47), .O(n451));
  andx g420(.A(n454), .B(n37), .O(n452));
  orx  g421(.A(pi02), .B(n44), .O(n453));
  invx g422(.A(n455), .O(n454));
  andx g423(.A(n457), .B(n456), .O(n455));
  orx  g424(.A(n459), .B(pi03), .O(n456));
  orx  g425(.A(n46), .B(n458), .O(n457));
  invx g426(.A(n459), .O(n458));
  orx  g427(.A(n461), .B(n460), .O(n459));
  andx g428(.A(n473), .B(po04), .O(n460));
  andx g429(.A(pi04), .B(n462), .O(n461));
  orx  g430(.A(n505), .B(n45), .O(n462));
  invx g431(.A(n464), .O(n463));
  orx  g432(.A(n466), .B(n465), .O(n464));
  andx g433(.A(n468), .B(n40), .O(n465));
  andx g434(.A(n467), .B(pi05), .O(n466));
  invx g435(.A(n468), .O(n467));
  orx  g436(.A(n474), .B(n469), .O(n468));
  andx g437(.A(n470), .B(po04), .O(n469));
  andx g438(.A(n472), .B(n471), .O(n470));
  orx  g439(.A(n36), .B(n557), .O(n471));
  orx  g440(.A(n473), .B(n558), .O(n472));
  invx g441(.A(n36), .O(n473));
  andx g442(.A(n562), .B(n505), .O(n474));
  invx g443(.A(n476), .O(n475));
  orx  g444(.A(n478), .B(n477), .O(n476));
  andx g445(.A(n480), .B(n540), .O(n477));
  andx g446(.A(n479), .B(pi07), .O(n478));
  invx g447(.A(n480), .O(n479));
  orx  g448(.A(n482), .B(n481), .O(n480));
  andx g449(.A(n571), .B(n505), .O(n481));
  andx g450(.A(n483), .B(po04), .O(n482));
  orx  g451(.A(n485), .B(n484), .O(n483));
  andx g452(.A(n567), .B(n553), .O(n484));
  invx g453(.A(n486), .O(n485));
  orx  g454(.A(n553), .B(n567), .O(n486));
  invx g455(.A(n488), .O(n487));
  orx  g456(.A(n490), .B(n489), .O(n488));
  andx g457(.A(n492), .B(n523), .O(n489));
  andx g458(.A(n491), .B(pi09), .O(n490));
  invx g459(.A(n492), .O(n491));
  orx  g460(.A(n497), .B(n493), .O(n492));
  andx g461(.A(n494), .B(po04), .O(n493));
  andx g462(.A(n496), .B(n495), .O(n494));
  orx  g463(.A(n538), .B(n551), .O(n495));
  invx g464(.A(n537), .O(n496));
  andx g465(.A(n543), .B(n505), .O(n497));
  invx g466(.A(n499), .O(n498));
  orx  g467(.A(n501), .B(n500), .O(n499));
  andx g468(.A(n503), .B(n695), .O(n500));
  andx g469(.A(n502), .B(pi11), .O(n501));
  invx g470(.A(n503), .O(n502));
  orx  g471(.A(n506), .B(n504), .O(n503));
  andx g472(.A(n526), .B(n505), .O(n504));
  invx g473(.A(po04), .O(n505));
  andx g474(.A(n517), .B(po04), .O(n506));
  orx  g475(.A(n509), .B(n508), .O(n507));
  andx g476(.A(n691), .B(n515), .O(n508));
  andx g477(.A(n510), .B(n692), .O(n509));
  andx g478(.A(n514), .B(n511), .O(n510));
  orx  g479(.A(n512), .B(n522), .O(n511));
  andx g480(.A(n513), .B(n535), .O(n512));
  invx g481(.A(n521), .O(n513));
  orx  g482(.A(n515), .B(n695), .O(n514));
  andx g483(.A(n33), .B(n516), .O(n515));
  invx g484(.A(n623), .O(n516));
  orx  g485(.A(n519), .B(n518), .O(n517));
  andx g486(.A(n521), .B(n535), .O(n518));
  invx g487(.A(n520), .O(n519));
  orx  g488(.A(n535), .B(n521), .O(n520));
  orx  g489(.A(n524), .B(n522), .O(n521));
  andx g490(.A(n526), .B(n523), .O(n522));
  invx g491(.A(pi09), .O(n523));
  andx g492(.A(n525), .B(pi09), .O(n524));
  invx g493(.A(n526), .O(n525));
  orx  g494(.A(n534), .B(n527), .O(n526));
  andx g495(.A(n528), .B(po06), .O(n527));
  andx g496(.A(n530), .B(n529), .O(n528));
  orx  g497(.A(n588), .B(n532), .O(n529));
  invx g498(.A(n531), .O(n530));
  andx g499(.A(n532), .B(n588), .O(n531));
  orx  g500(.A(n612), .B(n533), .O(n532));
  andx g501(.A(n42), .B(n615), .O(n533));
  andx g502(.A(n615), .B(n33), .O(n534));
  orx  g503(.A(n537), .B(n536), .O(n535));
  andx g504(.A(n543), .B(n540), .O(n536));
  andx g505(.A(n551), .B(n538), .O(n537));
  orx  g506(.A(n542), .B(n539), .O(n538));
  andx g507(.A(n541), .B(n540), .O(n539));
  invx g508(.A(pi07), .O(n540));
  invx g509(.A(n543), .O(n541));
  andx g510(.A(pi07), .B(n543), .O(n542));
  orx  g511(.A(n547), .B(n544), .O(n543));
  andx g512(.A(n600), .B(n545), .O(n544));
  orx  g513(.A(n546), .B(n33), .O(n545));
  andx g514(.A(n549), .B(n41), .O(n546));
  andx g515(.A(n548), .B(po06), .O(n547));
  andx g516(.A(n549), .B(n589), .O(n548));
  orx  g517(.A(n550), .B(n591), .O(n549));
  andx g518(.A(n598), .B(n597), .O(n550));
  orx  g519(.A(n552), .B(n568), .O(n551));
  andx g520(.A(n566), .B(n553), .O(n552));
  orx  g521(.A(n555), .B(n554), .O(n553));
  andx g522(.A(n562), .B(n46), .O(n554));
  andx g523(.A(n557), .B(n36), .O(n555));
  orx  g524(.A(pi04), .B(n701), .O(n556));
  invx g525(.A(n558), .O(n557));
  andx g526(.A(n560), .B(n559), .O(n558));
  orx  g527(.A(n562), .B(pi03), .O(n559));
  orx  g528(.A(n48), .B(n561), .O(n560));
  invx g529(.A(n562), .O(n561));
  orx  g530(.A(n564), .B(n563), .O(n562));
  andx g531(.A(po06), .B(n577), .O(n563));
  andx g532(.A(pi06), .B(n565), .O(n564));
  orx  g533(.A(n45), .B(n33), .O(n565));
  invx g534(.A(n567), .O(n566));
  orx  g535(.A(n569), .B(n568), .O(n567));
  andx g536(.A(n571), .B(n40), .O(n568));
  andx g537(.A(n570), .B(pi05), .O(n569));
  invx g538(.A(n571), .O(n570));
  orx  g539(.A(n580), .B(n572), .O(n571));
  andx g540(.A(n574), .B(n573), .O(n572));
  invx g541(.A(n593), .O(n573));
  andx g542(.A(po06), .B(n575), .O(n574));
  orx  g543(.A(n578), .B(n576), .O(n575));
  andx g544(.A(n577), .B(n48), .O(n576));
  invx g545(.A(n700), .O(n577));
  andx g546(.A(pi03), .B(n700), .O(n578));
  invx g547(.A(n33), .O(po06));
  andx g548(.A(n581), .B(n593), .O(n580));
  orx  g549(.A(n696), .B(n33), .O(n581));
  orx  g550(.A(n583), .B(n690), .O(n582));
  andx g551(.A(n622), .B(n584), .O(n583));
  orx  g552(.A(n586), .B(n585), .O(n584));
  andx g553(.A(pi09), .B(n623), .O(n585));
  andx g554(.A(n613), .B(n587), .O(n586));
  orx  g555(.A(n612), .B(n588), .O(n587));
  andx g556(.A(n598), .B(n589), .O(n588));
  invx g557(.A(n590), .O(n589));
  andx g558(.A(n597), .B(n591), .O(n590));
  orx  g559(.A(n592), .B(n699), .O(n591));
  andx g560(.A(n593), .B(n698), .O(n592));
  orx  g561(.A(n595), .B(n594), .O(n593));
  andx g562(.A(po08), .B(n606), .O(n594));
  andx g563(.A(pi08), .B(n596), .O(n595));
  orx  g564(.A(n44), .B(n625), .O(n596));
  orx  g565(.A(n40), .B(n600), .O(n597));
  orx  g566(.A(pi05), .B(n599), .O(n598));
  invx g567(.A(n600), .O(n599));
  orx  g568(.A(n608), .B(n601), .O(n600));
  andx g569(.A(n603), .B(n602), .O(n601));
  invx g570(.A(n645), .O(n602));
  andx g571(.A(po08), .B(n604), .O(n603));
  orx  g572(.A(n607), .B(n605), .O(n604));
  andx g573(.A(n606), .B(n47), .O(n605));
  invx g574(.A(n651), .O(n606));
  andx g575(.A(pi03), .B(n651), .O(n607));
  andx g576(.A(n609), .B(n645), .O(n608));
  orx  g577(.A(n610), .B(n625), .O(n609));
  orx  g578(.A(n643), .B(n611), .O(n610));
  invx g579(.A(n650), .O(n611));
  andx g580(.A(pi07), .B(n614), .O(n612));
  orx  g581(.A(pi07), .B(n614), .O(n613));
  invx g582(.A(n615), .O(n614));
  orx  g583(.A(n617), .B(n616), .O(n615));
  andx g584(.A(n634), .B(n625), .O(n616));
  andx g585(.A(n620), .B(n618), .O(n617));
  orx  g586(.A(n619), .B(n642), .O(n618));
  andx g587(.A(n629), .B(n633), .O(n619));
  orx  g588(.A(n621), .B(n630), .O(n620));
  andx g589(.A(po08), .B(n631), .O(n621));
  orx  g590(.A(pi09), .B(n623), .O(n622));
  orx  g591(.A(po08), .B(n654), .O(n623));
  invx g592(.A(n625), .O(po08));
  orx  g593(.A(n626), .B(n689), .O(n625));
  andx g594(.A(n653), .B(n627), .O(n626));
  orx  g595(.A(n652), .B(n628), .O(n627));
  andx g596(.A(n631), .B(n629), .O(n628));
  invx g597(.A(n630), .O(n629));
  andx g598(.A(n41), .B(n634), .O(n630));
  invx g599(.A(n632), .O(n631));
  andx g600(.A(n642), .B(n633), .O(n632));
  orx  g601(.A(n634), .B(n41), .O(n633));
  orx  g602(.A(n637), .B(n635), .O(n634));
  invx g603(.A(n636), .O(n635));
  orx  g604(.A(n638), .B(n668), .O(n636));
  andx g605(.A(n638), .B(n668), .O(n637));
  orx  g606(.A(n639), .B(n657), .O(n638));
  andx g607(.A(n641), .B(n640), .O(n639));
  orx  g608(.A(n647), .B(n47), .O(n640));
  orx  g609(.A(pi03), .B(n667), .O(n641));
  orx  g610(.A(n644), .B(n643), .O(n642));
  andx g611(.A(n46), .B(n651), .O(n643));
  andx g612(.A(n650), .B(n645), .O(n644));
  orx  g613(.A(n648), .B(n646), .O(n645));
  andx g614(.A(po10), .B(n647), .O(n646));
  invx g615(.A(n667), .O(n647));
  andx g616(.A(pi10), .B(n649), .O(n648));
  orx  g617(.A(n45), .B(n657), .O(n649));
  orx  g618(.A(n47), .B(n651), .O(n650));
  orx  g619(.A(pi08), .B(n44), .O(n651));
  andx g620(.A(pi07), .B(n654), .O(n652));
  orx  g621(.A(n654), .B(pi07), .O(n653));
  andx g622(.A(n661), .B(n655), .O(n654));
  orx  g623(.A(n671), .B(po10), .O(n655));
  invx g624(.A(n657), .O(po10));
  orx  g625(.A(n658), .B(n688), .O(n657));
  andx g626(.A(n659), .B(n670), .O(n658));
  orx  g627(.A(n660), .B(n662), .O(n659));
  andx g628(.A(pi05), .B(n671), .O(n660));
  orx  g629(.A(n670), .B(n662), .O(n661));
  invx g630(.A(n663), .O(n662));
  orx  g631(.A(n665), .B(n664), .O(n663));
  andx g632(.A(n667), .B(n668), .O(n664));
  andx g633(.A(n666), .B(n46), .O(n665));
  orx  g634(.A(n668), .B(n667), .O(n666));
  orx  g635(.A(pi10), .B(n45), .O(n667));
  andx g636(.A(n669), .B(pi12), .O(n668));
  orx  g637(.A(n674), .B(n701), .O(n669));
  orx  g638(.A(pi05), .B(n671), .O(n670));
  orx  g639(.A(n672), .B(n679), .O(n671));
  andx g640(.A(po12), .B(pi03), .O(n672));
  invx g641(.A(n674), .O(po12));
  orx  g642(.A(n688), .B(n675), .O(n674));
  orx  g643(.A(pi05), .B(n676), .O(n675));
  andx g644(.A(n678), .B(n677), .O(n676));
  orx  g645(.A(pi03), .B(n686), .O(n677));
  orx  g646(.A(n686), .B(n679), .O(n678));
  orx  g647(.A(n681), .B(n680), .O(n679));
  invx g648(.A(pi14), .O(n680));
  andx g649(.A(n684), .B(n682), .O(n681));
  andx g650(.A(n48), .B(n41), .O(n682));
  invx g651(.A(pi05), .O(n683));
  andx g652(.A(n685), .B(pi01), .O(n684));
  invx g653(.A(n688), .O(n685));
  andx g654(.A(n687), .B(pi01), .O(n686));
  invx g655(.A(pi12), .O(n687));
  orx  g656(.A(pi07), .B(n689), .O(n688));
  orx  g657(.A(pi09), .B(n690), .O(n689));
  invx g658(.A(n691), .O(n690));
  andx g659(.A(n695), .B(n692), .O(n691));
  andx g660(.A(n694), .B(n693), .O(n692));
  invx g661(.A(pi13), .O(n693));
  invx g662(.A(pi15), .O(n694));
  invx g663(.A(pi11), .O(n695));
  orx  g664(.A(n699), .B(n697), .O(n696));
  invx g665(.A(n698), .O(n697));
  orx  g666(.A(n46), .B(n700), .O(n698));
  andx g667(.A(n47), .B(n700), .O(n699));
  orx  g668(.A(pi06), .B(n44), .O(n700));
  invx g669(.A(pi01), .O(n701));
  invx g670(.A(pi03), .O(n702));
endmodule


