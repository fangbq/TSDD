// Benchmark "top" written by ABC on Fri Feb  7 13:28:40 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n510, n511, n512, n513, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
    n549, n550, n551, n552, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
    n588, n589, n590, n591, n593, n594, n595, n596, n598, n599, n600, n601,
    n603, n604, n605, n606, n608, n609, n610, n611, n613, n614, n615, n616,
    n618, n619, n620, n621, n622, n623, n624, n625, n627, n628, n629, n630,
    n632, n633, n634, n635, n637, n638, n639, n640, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n653, n654, n655, n656, n658, n659,
    n660, n661, n663, n664, n665, n666, n668, n669, n670, n671, n673, n674,
    n675, n676, n678, n679, n680, n681, n683, n684, n685, n686, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n699, n700, n701, n702,
    n704, n705, n706, n707, n709, n710, n711, n712, n714, n715, n716, n717,
    n719, n720, n721, n722, n724, n725, n726, n727;
  orx  g000(.a(pi30), .b(pi20), .O(n73));
  invx g001(.a(pi20), .O(n74));
  invx g002(.a(pi30), .O(n75));
  orx  g003(.a(n75), .b(n74), .O(n76));
  andx g004(.a(n76), .b(n73), .O(n77));
  invx g005(.a(pi12), .O(n78));
  orx  g006(.a(pi16), .b(n78), .O(n79));
  invx g007(.a(pi16), .O(n80));
  orx  g008(.a(n80), .b(pi12), .O(n81));
  andx g009(.a(n81), .b(n79), .O(n82));
  andx g010(.a(n82), .b(n77), .O(n83));
  andx g011(.a(n75), .b(n74), .O(n84));
  andx g012(.a(pi30), .b(pi20), .O(n85));
  orx  g013(.a(n85), .b(n84), .O(n86));
  andx g014(.a(n80), .b(pi12), .O(n87));
  andx g015(.a(pi16), .b(n78), .O(n88));
  orx  g016(.a(n88), .b(n87), .O(n89));
  andx g017(.a(n89), .b(n86), .O(n90));
  orx  g018(.a(n90), .b(n83), .O(n91));
  andx g019(.a(pi10), .b(pi01), .O(n92));
  invx g020(.a(pi07), .O(n93));
  invx g021(.a(pi32), .O(n94));
  andx g022(.a(n94), .b(n93), .O(n95));
  andx g023(.a(pi32), .b(pi07), .O(n96));
  orx  g024(.a(n96), .b(n95), .O(n97));
  invx g025(.a(pi17), .O(n98));
  andx g026(.a(n98), .b(pi08), .O(n99));
  invx g027(.a(pi08), .O(n100));
  andx g028(.a(pi17), .b(n100), .O(n101));
  orx  g029(.a(n101), .b(n99), .O(n102));
  orx  g030(.a(n102), .b(n97), .O(n103));
  orx  g031(.a(pi32), .b(pi07), .O(n104));
  orx  g032(.a(n94), .b(n93), .O(n105));
  andx g033(.a(n105), .b(n104), .O(n106));
  orx  g034(.a(pi17), .b(n100), .O(n107));
  orx  g035(.a(n98), .b(pi08), .O(n108));
  andx g036(.a(n108), .b(n107), .O(n109));
  orx  g037(.a(n109), .b(n106), .O(n110));
  andx g038(.a(n110), .b(n103), .O(n111));
  andx g039(.a(n111), .b(n92), .O(n112));
  invx g040(.a(n92), .O(n113));
  andx g041(.a(n109), .b(n106), .O(n114));
  andx g042(.a(n102), .b(n97), .O(n115));
  orx  g043(.a(n115), .b(n114), .O(n116));
  andx g044(.a(n116), .b(n113), .O(n117));
  orx  g045(.a(n117), .b(n112), .O(n118));
  orx  g046(.a(n118), .b(n91), .O(n119));
  orx  g047(.a(n89), .b(n86), .O(n120));
  orx  g048(.a(n82), .b(n77), .O(n121));
  andx g049(.a(n121), .b(n120), .O(n122));
  orx  g050(.a(n116), .b(n113), .O(n123));
  orx  g051(.a(n111), .b(n92), .O(n124));
  andx g052(.a(n124), .b(n123), .O(n125));
  orx  g053(.a(n125), .b(n122), .O(n126));
  andx g054(.a(n126), .b(n119), .O(n127));
  orx  g055(.a(pi36), .b(pi21), .O(n128));
  andx g056(.a(pi36), .b(pi21), .O(n129));
  invx g057(.a(n129), .O(n130));
  andx g058(.a(n130), .b(n128), .O(n131));
  invx g059(.a(pi35), .O(n132));
  andx g060(.a(n132), .b(pi22), .O(n133));
  invx g061(.a(pi22), .O(n134));
  andx g062(.a(pi35), .b(n134), .O(n135));
  orx  g063(.a(n135), .b(n133), .O(n136));
  andx g064(.a(n136), .b(n131), .O(n137));
  invx g065(.a(n137), .O(n138));
  orx  g066(.a(n136), .b(n131), .O(n139));
  andx g067(.a(n139), .b(n138), .O(n140));
  andx g068(.a(n140), .b(n127), .O(n141));
  andx g069(.a(n125), .b(n122), .O(n142));
  andx g070(.a(n118), .b(n91), .O(n143));
  orx  g071(.a(n143), .b(n142), .O(n144));
  invx g072(.a(n140), .O(n145));
  andx g073(.a(n145), .b(n144), .O(n146));
  orx  g074(.a(n146), .b(n141), .O(n147));
  andx g075(.a(pi01), .b(pi02), .O(n148));
  invx g076(.a(n148), .O(n149));
  orx  g077(.a(pi19), .b(pi31), .O(n150));
  invx g078(.a(pi31), .O(n151));
  invx g079(.a(pi19), .O(n152));
  orx  g080(.a(n152), .b(n151), .O(n153));
  andx g081(.a(n153), .b(n150), .O(n154));
  invx g082(.a(pi11), .O(n155));
  orx  g083(.a(pi15), .b(n155), .O(n156));
  invx g084(.a(pi15), .O(n157));
  orx  g085(.a(n157), .b(pi11), .O(n158));
  andx g086(.a(n158), .b(n156), .O(n159));
  andx g087(.a(n159), .b(n154), .O(n160));
  andx g088(.a(n152), .b(n151), .O(n161));
  andx g089(.a(pi19), .b(pi31), .O(n162));
  orx  g090(.a(n162), .b(n161), .O(n163));
  andx g091(.a(n157), .b(pi11), .O(n164));
  andx g092(.a(pi15), .b(n155), .O(n165));
  orx  g093(.a(n165), .b(n164), .O(n166));
  andx g094(.a(n166), .b(n163), .O(n167));
  orx  g095(.a(n167), .b(n160), .O(n168));
  orx  g096(.a(n168), .b(n149), .O(n169));
  orx  g097(.a(n166), .b(n163), .O(n170));
  orx  g098(.a(n159), .b(n154), .O(n171));
  andx g099(.a(n171), .b(n170), .O(n172));
  orx  g100(.a(n172), .b(n148), .O(n173));
  andx g101(.a(n173), .b(n169), .O(n174));
  invx g102(.a(pi05), .O(n175));
  invx g103(.a(pi29), .O(n176));
  andx g104(.a(n176), .b(n175), .O(n177));
  andx g105(.a(pi29), .b(pi05), .O(n178));
  orx  g106(.a(n178), .b(n177), .O(n179));
  invx g107(.a(pi18), .O(n180));
  andx g108(.a(n180), .b(pi06), .O(n181));
  invx g109(.a(pi06), .O(n182));
  andx g110(.a(pi18), .b(n182), .O(n183));
  orx  g111(.a(n183), .b(n181), .O(n184));
  orx  g112(.a(n184), .b(n179), .O(n185));
  andx g113(.a(n184), .b(n179), .O(n186));
  invx g114(.a(n186), .O(n187));
  andx g115(.a(n187), .b(n185), .O(n188));
  andx g116(.a(n188), .b(n174), .O(n189));
  andx g117(.a(n172), .b(n148), .O(n190));
  andx g118(.a(n168), .b(n149), .O(n191));
  orx  g119(.a(n191), .b(n190), .O(n192));
  invx g120(.a(n185), .O(n193));
  orx  g121(.a(n186), .b(n193), .O(n194));
  andx g122(.a(n194), .b(n192), .O(n195));
  orx  g123(.a(n195), .b(n189), .O(n196));
  orx  g124(.a(pi37), .b(pi26), .O(n197));
  andx g125(.a(pi37), .b(pi26), .O(n198));
  invx g126(.a(n198), .O(n199));
  andx g127(.a(n199), .b(n197), .O(n200));
  invx g128(.a(pi38), .O(n201));
  andx g129(.a(n201), .b(pi25), .O(n202));
  invx g130(.a(pi25), .O(n203));
  andx g131(.a(pi38), .b(n203), .O(n204));
  orx  g132(.a(n204), .b(n202), .O(n205));
  andx g133(.a(n205), .b(n200), .O(n206));
  invx g134(.a(n206), .O(n207));
  orx  g135(.a(n205), .b(n200), .O(n208));
  andx g136(.a(n208), .b(n207), .O(n209));
  invx g137(.a(n209), .O(n210));
  orx  g138(.a(n210), .b(n196), .O(n211));
  orx  g139(.a(n194), .b(n192), .O(n212));
  orx  g140(.a(n188), .b(n174), .O(n213));
  andx g141(.a(n213), .b(n212), .O(n214));
  orx  g142(.a(n209), .b(n214), .O(n215));
  andx g143(.a(n215), .b(n211), .O(n216));
  andx g144(.a(pi01), .b(pi03), .O(n217));
  invx g145(.a(n217), .O(n218));
  orx  g146(.a(n218), .b(n91), .O(n219));
  orx  g147(.a(n217), .b(n122), .O(n220));
  andx g148(.a(n220), .b(n219), .O(n221));
  andx g149(.a(n221), .b(n188), .O(n222));
  andx g150(.a(n217), .b(n122), .O(n223));
  andx g151(.a(n218), .b(n91), .O(n224));
  orx  g152(.a(n224), .b(n223), .O(n225));
  andx g153(.a(n225), .b(n194), .O(n226));
  orx  g154(.a(n226), .b(n222), .O(n227));
  orx  g155(.a(pi39), .b(pi28), .O(n228));
  andx g156(.a(pi39), .b(pi28), .O(n229));
  invx g157(.a(n229), .O(n230));
  andx g158(.a(n230), .b(n228), .O(n231));
  invx g159(.a(pi27), .O(n232));
  andx g160(.a(n232), .b(pi40), .O(n233));
  invx g161(.a(pi40), .O(n234));
  andx g162(.a(pi27), .b(n234), .O(n235));
  orx  g163(.a(n235), .b(n233), .O(n236));
  andx g164(.a(n236), .b(n231), .O(n237));
  invx g165(.a(n237), .O(n238));
  orx  g166(.a(n236), .b(n231), .O(n239));
  andx g167(.a(n239), .b(n238), .O(n240));
  invx g168(.a(n240), .O(n241));
  orx  g169(.a(n241), .b(n227), .O(n242));
  orx  g170(.a(n225), .b(n194), .O(n243));
  orx  g171(.a(n221), .b(n188), .O(n244));
  andx g172(.a(n244), .b(n243), .O(n245));
  orx  g173(.a(n240), .b(n245), .O(n246));
  andx g174(.a(n246), .b(n242), .O(n247));
  orx  g175(.a(n247), .b(n216), .O(n248));
  andx g176(.a(pi01), .b(pi09), .O(n249));
  andx g177(.a(n249), .b(n111), .O(n250));
  invx g178(.a(n249), .O(n251));
  andx g179(.a(n251), .b(n116), .O(n252));
  orx  g180(.a(n252), .b(n250), .O(n253));
  orx  g181(.a(n253), .b(n168), .O(n254));
  orx  g182(.a(n251), .b(n116), .O(n255));
  orx  g183(.a(n249), .b(n111), .O(n256));
  andx g184(.a(n256), .b(n255), .O(n257));
  orx  g185(.a(n257), .b(n172), .O(n258));
  andx g186(.a(n258), .b(n254), .O(n259));
  orx  g187(.a(pi34), .b(pi23), .O(n260));
  andx g188(.a(pi34), .b(pi23), .O(n261));
  invx g189(.a(n261), .O(n262));
  andx g190(.a(n262), .b(n260), .O(n263));
  invx g191(.a(pi24), .O(n264));
  andx g192(.a(n264), .b(pi33), .O(n265));
  invx g193(.a(pi33), .O(n266));
  andx g194(.a(pi24), .b(n266), .O(n267));
  orx  g195(.a(n267), .b(n265), .O(n268));
  andx g196(.a(n268), .b(n263), .O(n269));
  invx g197(.a(n269), .O(n270));
  orx  g198(.a(n268), .b(n263), .O(n271));
  andx g199(.a(n271), .b(n270), .O(n272));
  andx g200(.a(n272), .b(n259), .O(n273));
  andx g201(.a(n257), .b(n172), .O(n274));
  andx g202(.a(n253), .b(n168), .O(n275));
  orx  g203(.a(n275), .b(n274), .O(n276));
  invx g204(.a(n272), .O(n277));
  andx g205(.a(n277), .b(n276), .O(n278));
  orx  g206(.a(n278), .b(n273), .O(n279));
  andx g207(.a(n279), .b(n147), .O(n280));
  orx  g208(.a(n145), .b(n144), .O(n281));
  orx  g209(.a(n140), .b(n127), .O(n282));
  andx g210(.a(n282), .b(n281), .O(n283));
  orx  g211(.a(n277), .b(n276), .O(n284));
  orx  g212(.a(n272), .b(n259), .O(n285));
  andx g213(.a(n285), .b(n284), .O(n286));
  andx g214(.a(n286), .b(n283), .O(n287));
  orx  g215(.a(n287), .b(n280), .O(n288));
  orx  g216(.a(n288), .b(n248), .O(n289));
  orx  g217(.a(n286), .b(n283), .O(n290));
  andx g218(.a(n209), .b(n214), .O(n291));
  andx g219(.a(n210), .b(n196), .O(n292));
  orx  g220(.a(n292), .b(n291), .O(n293));
  andx g221(.a(n240), .b(n245), .O(n294));
  andx g222(.a(n241), .b(n227), .O(n295));
  orx  g223(.a(n295), .b(n294), .O(n296));
  andx g224(.a(n296), .b(n293), .O(n297));
  andx g225(.a(n247), .b(n216), .O(n298));
  orx  g226(.a(n298), .b(n297), .O(n299));
  orx  g227(.a(n299), .b(n290), .O(n300));
  andx g228(.a(n300), .b(n289), .O(n301));
  andx g229(.a(pi01), .b(pi14), .O(n302));
  andx g230(.a(n203), .b(n134), .O(n303));
  andx g231(.a(pi25), .b(pi22), .O(n304));
  orx  g232(.a(n304), .b(n303), .O(n305));
  andx g233(.a(n266), .b(pi40), .O(n306));
  andx g234(.a(pi33), .b(n234), .O(n307));
  orx  g235(.a(n307), .b(n306), .O(n308));
  orx  g236(.a(n308), .b(n305), .O(n309));
  orx  g237(.a(pi25), .b(pi22), .O(n310));
  orx  g238(.a(n203), .b(n134), .O(n311));
  andx g239(.a(n311), .b(n310), .O(n312));
  orx  g240(.a(pi33), .b(n234), .O(n313));
  orx  g241(.a(n266), .b(pi40), .O(n314));
  andx g242(.a(n314), .b(n313), .O(n315));
  orx  g243(.a(n315), .b(n312), .O(n316));
  andx g244(.a(n316), .b(n309), .O(n317));
  andx g245(.a(n317), .b(n302), .O(n318));
  invx g246(.a(n302), .O(n319));
  andx g247(.a(n315), .b(n312), .O(n320));
  andx g248(.a(n308), .b(n305), .O(n321));
  orx  g249(.a(n321), .b(n320), .O(n322));
  andx g250(.a(n322), .b(n319), .O(n323));
  orx  g251(.a(n323), .b(n318), .O(n324));
  orx  g252(.a(pi26), .b(pi21), .O(n325));
  invx g253(.a(pi21), .O(n326));
  invx g254(.a(pi26), .O(n327));
  orx  g255(.a(n327), .b(n326), .O(n328));
  andx g256(.a(n328), .b(n325), .O(n329));
  invx g257(.a(pi34), .O(n330));
  orx  g258(.a(pi39), .b(n330), .O(n331));
  invx g259(.a(pi39), .O(n332));
  orx  g260(.a(n332), .b(pi34), .O(n333));
  andx g261(.a(n333), .b(n331), .O(n334));
  andx g262(.a(n334), .b(n329), .O(n335));
  andx g263(.a(n327), .b(n326), .O(n336));
  andx g264(.a(pi26), .b(pi21), .O(n337));
  orx  g265(.a(n337), .b(n336), .O(n338));
  andx g266(.a(n332), .b(pi34), .O(n339));
  andx g267(.a(pi39), .b(n330), .O(n340));
  orx  g268(.a(n340), .b(n339), .O(n341));
  andx g269(.a(n341), .b(n338), .O(n342));
  orx  g270(.a(n342), .b(n335), .O(n343));
  orx  g271(.a(n343), .b(n324), .O(n344));
  orx  g272(.a(n322), .b(n319), .O(n345));
  orx  g273(.a(n317), .b(n302), .O(n346));
  andx g274(.a(n346), .b(n345), .O(n347));
  orx  g275(.a(n341), .b(n338), .O(n348));
  orx  g276(.a(n334), .b(n329), .O(n349));
  andx g277(.a(n349), .b(n348), .O(n350));
  orx  g278(.a(n350), .b(n347), .O(n351));
  andx g279(.a(n351), .b(n344), .O(n352));
  orx  g280(.a(pi31), .b(pi32), .O(n353));
  andx g281(.a(pi31), .b(pi32), .O(n354));
  invx g282(.a(n354), .O(n355));
  andx g283(.a(n355), .b(n353), .O(n356));
  andx g284(.a(n75), .b(pi29), .O(n357));
  andx g285(.a(pi30), .b(n176), .O(n358));
  orx  g286(.a(n358), .b(n357), .O(n359));
  andx g287(.a(n359), .b(n356), .O(n360));
  invx g288(.a(n360), .O(n361));
  orx  g289(.a(n359), .b(n356), .O(n362));
  andx g290(.a(n362), .b(n361), .O(n363));
  andx g291(.a(n363), .b(n352), .O(n364));
  andx g292(.a(n350), .b(n347), .O(n365));
  andx g293(.a(n343), .b(n324), .O(n366));
  orx  g294(.a(n366), .b(n365), .O(n367));
  invx g295(.a(n363), .O(n368));
  andx g296(.a(n368), .b(n367), .O(n369));
  orx  g297(.a(n369), .b(n364), .O(n370));
  andx g298(.a(pi01), .b(pi13), .O(n371));
  andx g299(.a(n371), .b(n317), .O(n372));
  invx g300(.a(n371), .O(n373));
  andx g301(.a(n373), .b(n322), .O(n374));
  orx  g302(.a(n374), .b(n372), .O(n375));
  orx  g303(.a(pi38), .b(pi35), .O(n376));
  orx  g304(.a(n201), .b(n132), .O(n377));
  andx g305(.a(n377), .b(n376), .O(n378));
  orx  g306(.a(pi24), .b(n232), .O(n379));
  orx  g307(.a(n264), .b(pi27), .O(n380));
  andx g308(.a(n380), .b(n379), .O(n381));
  andx g309(.a(n381), .b(n378), .O(n382));
  andx g310(.a(n201), .b(n132), .O(n383));
  andx g311(.a(pi38), .b(pi35), .O(n384));
  orx  g312(.a(n384), .b(n383), .O(n385));
  andx g313(.a(n264), .b(pi27), .O(n386));
  andx g314(.a(pi24), .b(n232), .O(n387));
  orx  g315(.a(n387), .b(n386), .O(n388));
  andx g316(.a(n388), .b(n385), .O(n389));
  orx  g317(.a(n389), .b(n382), .O(n390));
  orx  g318(.a(n390), .b(n375), .O(n391));
  orx  g319(.a(n373), .b(n322), .O(n392));
  orx  g320(.a(n371), .b(n317), .O(n393));
  andx g321(.a(n393), .b(n392), .O(n394));
  orx  g322(.a(n388), .b(n385), .O(n395));
  orx  g323(.a(n381), .b(n378), .O(n396));
  andx g324(.a(n396), .b(n395), .O(n397));
  orx  g325(.a(n397), .b(n394), .O(n398));
  andx g326(.a(n398), .b(n391), .O(n399));
  orx  g327(.a(pi17), .b(pi15), .O(n400));
  andx g328(.a(pi17), .b(pi15), .O(n401));
  invx g329(.a(n401), .O(n402));
  andx g330(.a(n402), .b(n400), .O(n403));
  andx g331(.a(n80), .b(pi18), .O(n404));
  andx g332(.a(pi16), .b(n180), .O(n405));
  orx  g333(.a(n405), .b(n404), .O(n406));
  andx g334(.a(n406), .b(n403), .O(n407));
  invx g335(.a(n407), .O(n408));
  orx  g336(.a(n406), .b(n403), .O(n409));
  andx g337(.a(n409), .b(n408), .O(n410));
  andx g338(.a(n410), .b(n399), .O(n411));
  andx g339(.a(n397), .b(n394), .O(n412));
  andx g340(.a(n390), .b(n375), .O(n413));
  orx  g341(.a(n413), .b(n412), .O(n414));
  invx g342(.a(n410), .O(n415));
  andx g343(.a(n415), .b(n414), .O(n416));
  orx  g344(.a(n416), .b(n411), .O(n417));
  andx g345(.a(n417), .b(n370), .O(n418));
  andx g346(.a(pi01), .b(pi04), .O(n419));
  invx g347(.a(n419), .O(n420));
  orx  g348(.a(n420), .b(n343), .O(n421));
  orx  g349(.a(n419), .b(n350), .O(n422));
  andx g350(.a(n422), .b(n421), .O(n423));
  invx g351(.a(pi36), .O(n424));
  invx g352(.a(pi37), .O(n425));
  andx g353(.a(n425), .b(n424), .O(n426));
  andx g354(.a(pi37), .b(pi36), .O(n427));
  orx  g355(.a(n427), .b(n426), .O(n428));
  invx g356(.a(pi23), .O(n429));
  andx g357(.a(n429), .b(pi28), .O(n430));
  invx g358(.a(pi28), .O(n431));
  andx g359(.a(pi23), .b(n431), .O(n432));
  orx  g360(.a(n432), .b(n430), .O(n433));
  orx  g361(.a(n433), .b(n428), .O(n434));
  andx g362(.a(n433), .b(n428), .O(n435));
  invx g363(.a(n435), .O(n436));
  andx g364(.a(n436), .b(n434), .O(n437));
  andx g365(.a(n437), .b(n423), .O(n438));
  andx g366(.a(n419), .b(n350), .O(n439));
  andx g367(.a(n420), .b(n343), .O(n440));
  orx  g368(.a(n440), .b(n439), .O(n441));
  invx g369(.a(n434), .O(n442));
  orx  g370(.a(n435), .b(n442), .O(n443));
  andx g371(.a(n443), .b(n441), .O(n444));
  orx  g372(.a(n444), .b(n438), .O(n445));
  orx  g373(.a(pi08), .b(pi11), .O(n446));
  andx g374(.a(pi08), .b(pi11), .O(n447));
  invx g375(.a(n447), .O(n448));
  andx g376(.a(n448), .b(n446), .O(n449));
  andx g377(.a(n78), .b(pi06), .O(n450));
  andx g378(.a(pi12), .b(n182), .O(n451));
  orx  g379(.a(n451), .b(n450), .O(n452));
  andx g380(.a(n452), .b(n449), .O(n453));
  invx g381(.a(n453), .O(n454));
  orx  g382(.a(n452), .b(n449), .O(n455));
  andx g383(.a(n455), .b(n454), .O(n456));
  invx g384(.a(n456), .O(n457));
  orx  g385(.a(n457), .b(n445), .O(n458));
  orx  g386(.a(n443), .b(n441), .O(n459));
  orx  g387(.a(n437), .b(n423), .O(n460));
  andx g388(.a(n460), .b(n459), .O(n461));
  orx  g389(.a(n456), .b(n461), .O(n462));
  andx g390(.a(n462), .b(n458), .O(n463));
  andx g391(.a(pi01), .b(pi00), .O(n464));
  invx g392(.a(n464), .O(n465));
  orx  g393(.a(n465), .b(n390), .O(n466));
  orx  g394(.a(n464), .b(n397), .O(n467));
  andx g395(.a(n467), .b(n466), .O(n468));
  andx g396(.a(n468), .b(n437), .O(n469));
  andx g397(.a(n464), .b(n397), .O(n470));
  andx g398(.a(n465), .b(n390), .O(n471));
  orx  g399(.a(n471), .b(n470), .O(n472));
  andx g400(.a(n472), .b(n443), .O(n473));
  orx  g401(.a(n473), .b(n469), .O(n474));
  orx  g402(.a(pi19), .b(pi07), .O(n475));
  andx g403(.a(pi19), .b(pi07), .O(n476));
  invx g404(.a(n476), .O(n477));
  andx g405(.a(n477), .b(n475), .O(n478));
  andx g406(.a(n74), .b(pi05), .O(n479));
  andx g407(.a(pi20), .b(n175), .O(n480));
  orx  g408(.a(n480), .b(n479), .O(n481));
  andx g409(.a(n481), .b(n478), .O(n482));
  invx g410(.a(n482), .O(n483));
  orx  g411(.a(n481), .b(n478), .O(n484));
  andx g412(.a(n484), .b(n483), .O(n485));
  invx g413(.a(n485), .O(n486));
  orx  g414(.a(n486), .b(n474), .O(n487));
  orx  g415(.a(n472), .b(n443), .O(n488));
  orx  g416(.a(n468), .b(n437), .O(n489));
  andx g417(.a(n489), .b(n488), .O(n490));
  orx  g418(.a(n485), .b(n490), .O(n491));
  andx g419(.a(n491), .b(n487), .O(n492));
  andx g420(.a(n492), .b(n463), .O(n493));
  andx g421(.a(n493), .b(n418), .O(n494));
  invx g422(.a(n494), .O(n495));
  orx  g423(.a(n495), .b(n301), .O(n496));
  orx  g424(.a(n496), .b(n147), .O(n497));
  andx g425(.a(n497), .b(pi36), .O(n498));
  orx  g426(.a(n279), .b(n147), .O(n499));
  andx g427(.a(n499), .b(n290), .O(n500));
  andx g428(.a(n500), .b(n297), .O(n501));
  orx  g429(.a(n296), .b(n293), .O(n502));
  andx g430(.a(n502), .b(n248), .O(n503));
  andx g431(.a(n503), .b(n280), .O(n504));
  orx  g432(.a(n504), .b(n501), .O(n505));
  andx g433(.a(n494), .b(n505), .O(n506));
  andx g434(.a(n506), .b(n283), .O(n507));
  andx g435(.a(n507), .b(n424), .O(n508));
  orx  g436(.a(n508), .b(n498), .O(po00));
  orx  g437(.a(n496), .b(n293), .O(n510));
  andx g438(.a(n510), .b(pi37), .O(n511));
  andx g439(.a(n506), .b(n216), .O(n512));
  andx g440(.a(n512), .b(n425), .O(n513));
  orx  g441(.a(n513), .b(n511), .O(po01));
  andx g442(.a(n485), .b(n490), .O(n515));
  andx g443(.a(n486), .b(n474), .O(n516));
  orx  g444(.a(n516), .b(n515), .O(n517));
  andx g445(.a(n517), .b(n463), .O(n518));
  orx  g446(.a(n368), .b(n367), .O(n519));
  orx  g447(.a(n363), .b(n352), .O(n520));
  andx g448(.a(n520), .b(n519), .O(n521));
  andx g449(.a(n417), .b(n521), .O(n522));
  andx g450(.a(n522), .b(n518), .O(n523));
  invx g451(.a(n523), .O(n524));
  orx  g452(.a(n524), .b(n301), .O(n525));
  orx  g453(.a(n525), .b(n296), .O(n526));
  andx g454(.a(n526), .b(pi39), .O(n527));
  andx g455(.a(n523), .b(n505), .O(n528));
  andx g456(.a(n528), .b(n247), .O(n529));
  andx g457(.a(n529), .b(n332), .O(n530));
  orx  g458(.a(n530), .b(n527), .O(po02));
  orx  g459(.a(n415), .b(n414), .O(n532));
  orx  g460(.a(n410), .b(n399), .O(n533));
  andx g461(.a(n533), .b(n532), .O(n534));
  andx g462(.a(n534), .b(n521), .O(n535));
  andx g463(.a(n456), .b(n461), .O(n536));
  andx g464(.a(n457), .b(n445), .O(n537));
  orx  g465(.a(n537), .b(n536), .O(n538));
  andx g466(.a(n517), .b(n538), .O(n539));
  andx g467(.a(n539), .b(n535), .O(n540));
  invx g468(.a(n540), .O(n541));
  orx  g469(.a(n541), .b(n301), .O(n542));
  orx  g470(.a(n542), .b(n296), .O(n543));
  andx g471(.a(n543), .b(pi40), .O(n544));
  andx g472(.a(n540), .b(n505), .O(n545));
  andx g473(.a(n545), .b(n247), .O(n546));
  andx g474(.a(n546), .b(n234), .O(n547));
  orx  g475(.a(n547), .b(n544), .O(po03));
  orx  g476(.a(n496), .b(n296), .O(n549));
  andx g477(.a(n549), .b(pi28), .O(n550));
  andx g478(.a(n506), .b(n247), .O(n551));
  andx g479(.a(n551), .b(n431), .O(n552));
  orx  g480(.a(n552), .b(n550), .O(po04));
  andx g481(.a(n538), .b(n534), .O(n554));
  andx g482(.a(n492), .b(n370), .O(n555));
  andx g483(.a(n555), .b(n554), .O(n556));
  invx g484(.a(n556), .O(n557));
  orx  g485(.a(n557), .b(n301), .O(n558));
  orx  g486(.a(n558), .b(n279), .O(n559));
  andx g487(.a(n559), .b(pi24), .O(n560));
  andx g488(.a(n556), .b(n505), .O(n561));
  andx g489(.a(n561), .b(n286), .O(n562));
  andx g490(.a(n562), .b(n264), .O(n563));
  orx  g491(.a(n563), .b(n560), .O(po05));
  orx  g492(.a(n534), .b(n521), .O(n565));
  orx  g493(.a(n539), .b(n493), .O(n566));
  orx  g494(.a(n566), .b(n565), .O(n567));
  orx  g495(.a(n492), .b(n463), .O(n568));
  orx  g496(.a(n568), .b(n418), .O(n569));
  orx  g497(.a(n569), .b(n535), .O(n570));
  andx g498(.a(n570), .b(n567), .O(n571));
  andx g499(.a(n298), .b(n280), .O(n572));
  invx g500(.a(n572), .O(n573));
  orx  g501(.a(n573), .b(n571), .O(n574));
  orx  g502(.a(n574), .b(n417), .O(n575));
  andx g503(.a(n575), .b(pi18), .O(n576));
  orx  g504(.a(n517), .b(n538), .O(n577));
  andx g505(.a(n568), .b(n577), .O(n578));
  andx g506(.a(n578), .b(n418), .O(n579));
  orx  g507(.a(n417), .b(n370), .O(n580));
  andx g508(.a(n539), .b(n565), .O(n581));
  andx g509(.a(n581), .b(n580), .O(n582));
  orx  g510(.a(n582), .b(n579), .O(n583));
  andx g511(.a(n572), .b(n583), .O(n584));
  andx g512(.a(n584), .b(n534), .O(n585));
  andx g513(.a(n585), .b(n180), .O(n586));
  orx  g514(.a(n586), .b(n576), .O(po06));
  orx  g515(.a(n574), .b(n538), .O(n588));
  andx g516(.a(n588), .b(pi06), .O(n589));
  andx g517(.a(n584), .b(n463), .O(n590));
  andx g518(.a(n590), .b(n182), .O(n591));
  orx  g519(.a(n591), .b(n589), .O(po07));
  orx  g520(.a(n574), .b(n517), .O(n593));
  andx g521(.a(n593), .b(pi05), .O(n594));
  andx g522(.a(n584), .b(n492), .O(n595));
  andx g523(.a(n595), .b(n175), .O(n596));
  orx  g524(.a(n596), .b(n594), .O(po08));
  orx  g525(.a(n542), .b(n279), .O(n598));
  andx g526(.a(n598), .b(pi33), .O(n599));
  andx g527(.a(n545), .b(n286), .O(n600));
  andx g528(.a(n600), .b(n266), .O(n601));
  orx  g529(.a(n601), .b(n599), .O(po09));
  orx  g530(.a(n496), .b(n279), .O(n603));
  andx g531(.a(n603), .b(pi23), .O(n604));
  andx g532(.a(n506), .b(n286), .O(n605));
  andx g533(.a(n605), .b(n429), .O(n606));
  orx  g534(.a(n606), .b(n604), .O(po10));
  orx  g535(.a(n558), .b(n147), .O(n608));
  andx g536(.a(n608), .b(pi35), .O(n609));
  andx g537(.a(n561), .b(n283), .O(n610));
  andx g538(.a(n610), .b(n132), .O(n611));
  orx  g539(.a(n611), .b(n609), .O(po11));
  orx  g540(.a(n574), .b(n370), .O(n613));
  andx g541(.a(n613), .b(pi29), .O(n614));
  andx g542(.a(n584), .b(n521), .O(n615));
  andx g543(.a(n615), .b(n176), .O(n616));
  orx  g544(.a(n616), .b(n614), .O(po12));
  andx g545(.a(n287), .b(n297), .O(n618));
  invx g546(.a(n618), .O(n619));
  orx  g547(.a(n619), .b(n571), .O(n620));
  orx  g548(.a(n620), .b(n417), .O(n621));
  andx g549(.a(n621), .b(pi17), .O(n622));
  andx g550(.a(n618), .b(n583), .O(n623));
  andx g551(.a(n623), .b(n534), .O(n624));
  andx g552(.a(n624), .b(n98), .O(n625));
  orx  g553(.a(n625), .b(n622), .O(po13));
  orx  g554(.a(n620), .b(n538), .O(n627));
  andx g555(.a(n627), .b(pi08), .O(n628));
  andx g556(.a(n623), .b(n463), .O(n629));
  andx g557(.a(n629), .b(n100), .O(n630));
  orx  g558(.a(n630), .b(n628), .O(po14));
  orx  g559(.a(n620), .b(n517), .O(n632));
  andx g560(.a(n632), .b(pi07), .O(n633));
  andx g561(.a(n623), .b(n492), .O(n634));
  andx g562(.a(n634), .b(n93), .O(n635));
  orx  g563(.a(n635), .b(n633), .O(po15));
  orx  g564(.a(n620), .b(n370), .O(n637));
  andx g565(.a(n637), .b(pi32), .O(n638));
  andx g566(.a(n623), .b(n521), .O(n639));
  andx g567(.a(n639), .b(n94), .O(n640));
  orx  g568(.a(n640), .b(n638), .O(po16));
  andx g569(.a(n296), .b(n216), .O(n642));
  andx g570(.a(n286), .b(n147), .O(n643));
  andx g571(.a(n643), .b(n642), .O(n644));
  invx g572(.a(n644), .O(n645));
  orx  g573(.a(n645), .b(n571), .O(n646));
  orx  g574(.a(n646), .b(n417), .O(n647));
  andx g575(.a(n647), .b(pi15), .O(n648));
  andx g576(.a(n644), .b(n583), .O(n649));
  andx g577(.a(n649), .b(n534), .O(n650));
  andx g578(.a(n650), .b(n157), .O(n651));
  orx  g579(.a(n651), .b(n648), .O(po17));
  orx  g580(.a(n646), .b(n538), .O(n653));
  andx g581(.a(n653), .b(pi11), .O(n654));
  andx g582(.a(n649), .b(n463), .O(n655));
  andx g583(.a(n655), .b(n155), .O(n656));
  orx  g584(.a(n656), .b(n654), .O(po18));
  orx  g585(.a(n646), .b(n517), .O(n658));
  andx g586(.a(n658), .b(pi19), .O(n659));
  andx g587(.a(n649), .b(n492), .O(n660));
  andx g588(.a(n660), .b(n152), .O(n661));
  orx  g589(.a(n661), .b(n659), .O(po19));
  orx  g590(.a(n646), .b(n370), .O(n663));
  andx g591(.a(n663), .b(pi31), .O(n664));
  andx g592(.a(n649), .b(n521), .O(n665));
  andx g593(.a(n665), .b(n151), .O(n666));
  orx  g594(.a(n666), .b(n664), .O(po20));
  orx  g595(.a(n542), .b(n147), .O(n668));
  andx g596(.a(n668), .b(pi22), .O(n669));
  andx g597(.a(n545), .b(n283), .O(n670));
  andx g598(.a(n670), .b(n134), .O(n671));
  orx  g599(.a(n671), .b(n669), .O(po21));
  orx  g600(.a(n525), .b(n279), .O(n673));
  andx g601(.a(n673), .b(pi34), .O(n674));
  andx g602(.a(n528), .b(n286), .O(n675));
  andx g603(.a(n675), .b(n330), .O(n676));
  orx  g604(.a(n676), .b(n674), .O(po22));
  orx  g605(.a(n525), .b(n147), .O(n678));
  andx g606(.a(n678), .b(pi21), .O(n679));
  andx g607(.a(n528), .b(n283), .O(n680));
  andx g608(.a(n680), .b(n326), .O(n681));
  orx  g609(.a(n681), .b(n679), .O(po23));
  orx  g610(.a(n525), .b(n293), .O(n683));
  andx g611(.a(n683), .b(pi26), .O(n684));
  andx g612(.a(n528), .b(n216), .O(n685));
  andx g613(.a(n685), .b(n327), .O(n686));
  orx  g614(.a(n686), .b(n684), .O(po24));
  andx g615(.a(n247), .b(n293), .O(n688));
  andx g616(.a(n279), .b(n283), .O(n689));
  andx g617(.a(n689), .b(n688), .O(n690));
  invx g618(.a(n690), .O(n691));
  orx  g619(.a(n691), .b(n571), .O(n692));
  orx  g620(.a(n692), .b(n417), .O(n693));
  andx g621(.a(n693), .b(pi16), .O(n694));
  andx g622(.a(n690), .b(n583), .O(n695));
  andx g623(.a(n695), .b(n534), .O(n696));
  andx g624(.a(n696), .b(n80), .O(n697));
  orx  g625(.a(n697), .b(n694), .O(po25));
  orx  g626(.a(n692), .b(n538), .O(n699));
  andx g627(.a(n699), .b(pi12), .O(n700));
  andx g628(.a(n695), .b(n463), .O(n701));
  andx g629(.a(n701), .b(n78), .O(n702));
  orx  g630(.a(n702), .b(n700), .O(po26));
  orx  g631(.a(n692), .b(n517), .O(n704));
  andx g632(.a(n704), .b(pi20), .O(n705));
  andx g633(.a(n695), .b(n492), .O(n706));
  andx g634(.a(n706), .b(n74), .O(n707));
  orx  g635(.a(n707), .b(n705), .O(po27));
  orx  g636(.a(n692), .b(n370), .O(n709));
  andx g637(.a(n709), .b(pi30), .O(n710));
  andx g638(.a(n695), .b(n521), .O(n711));
  andx g639(.a(n711), .b(n75), .O(n712));
  orx  g640(.a(n712), .b(n710), .O(po28));
  orx  g641(.a(n558), .b(n293), .O(n714));
  andx g642(.a(n714), .b(pi38), .O(n715));
  andx g643(.a(n561), .b(n216), .O(n716));
  andx g644(.a(n716), .b(n201), .O(n717));
  orx  g645(.a(n717), .b(n715), .O(po29));
  orx  g646(.a(n542), .b(n293), .O(n719));
  andx g647(.a(n719), .b(pi25), .O(n720));
  andx g648(.a(n545), .b(n216), .O(n721));
  andx g649(.a(n721), .b(n203), .O(n722));
  orx  g650(.a(n722), .b(n720), .O(po30));
  orx  g651(.a(n558), .b(n296), .O(n724));
  andx g652(.a(n724), .b(pi27), .O(n725));
  andx g653(.a(n561), .b(n247), .O(n726));
  andx g654(.a(n726), .b(n232), .O(n727));
  orx  g655(.a(n727), .b(n725), .O(po31));
endmodule


