// Benchmark "unsigned_mult" written by ABC on Fri Feb  7 13:49:25 2014

module unsigned_mult ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19;
  wire n40, n41, n43, n44, n45, n46, n47, n49, n50, n51, n52, n53, n54, n55,
    n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69, n71, n72,
    n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n85, n86, n87, n88,
    n89, n91, n92, n93, n94, n95, n96, n97, n98, n100, n101, n102, n103,
    n104, n105, n107, n108, n109, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161;
  bufx g0000(.A(n1161), .O(n40));
  bufx g0001(.A(n1150), .O(n41));
  orx  g0002(.A(n44), .B(n43), .O(po09));
  andx g0003(.A(n807), .B(n46), .O(n43));
  invx g0004(.A(n45), .O(n44));
  orx  g0005(.A(n46), .B(n807), .O(n45));
  orx  g0006(.A(n716), .B(n47), .O(n46));
  invx g0007(.A(n718), .O(n47));
  andx g0008(.A(n50), .B(n49), .O(po08));
  orx  g0009(.A(n800), .B(n52), .O(n49));
  orx  g0010(.A(n51), .B(n799), .O(n50));
  invx g0011(.A(n52), .O(n51));
  orx  g0012(.A(n53), .B(n720), .O(n52));
  andx g0013(.A(n55), .B(n54), .O(n53));
  orx  g0014(.A(n105), .B(n895), .O(n54));
  invx g0015(.A(n723), .O(n55));
  orx  g0016(.A(n58), .B(n57), .O(po07));
  andx g0017(.A(n790), .B(n60), .O(n57));
  invx g0018(.A(n59), .O(n58));
  orx  g0019(.A(n60), .B(n790), .O(n59));
  orx  g0020(.A(n724), .B(n61), .O(n60));
  invx g0021(.A(n726), .O(n61));
  andx g0022(.A(n64), .B(n63), .O(po06));
  orx  g0023(.A(n783), .B(n66), .O(n63));
  orx  g0024(.A(n65), .B(n782), .O(n64));
  invx g0025(.A(n66), .O(n65));
  orx  g0026(.A(n67), .B(n728), .O(n66));
  andx g0027(.A(n69), .B(n68), .O(n67));
  orx  g0028(.A(n105), .B(n1031), .O(n68));
  invx g0029(.A(n731), .O(n69));
  orx  g0030(.A(n72), .B(n71), .O(po05));
  andx g0031(.A(n773), .B(n74), .O(n71));
  invx g0032(.A(n73), .O(n72));
  orx  g0033(.A(n74), .B(n773), .O(n73));
  orx  g0034(.A(n732), .B(n75), .O(n74));
  invx g0035(.A(n734), .O(n75));
  andx g0036(.A(n78), .B(n77), .O(po04));
  orx  g0037(.A(n766), .B(n80), .O(n77));
  orx  g0038(.A(n79), .B(n765), .O(n78));
  invx g0039(.A(n80), .O(n79));
  orx  g0040(.A(n81), .B(n736), .O(n80));
  andx g0041(.A(n83), .B(n82), .O(n81));
  orx  g0042(.A(n105), .B(n1117), .O(n82));
  invx g0043(.A(n739), .O(n83));
  orx  g0044(.A(n86), .B(n85), .O(po03));
  andx g0045(.A(n756), .B(n88), .O(n85));
  invx g0046(.A(n87), .O(n86));
  orx  g0047(.A(n88), .B(n756), .O(n87));
  orx  g0048(.A(n740), .B(n89), .O(n88));
  invx g0049(.A(n742), .O(n89));
  orx  g0050(.A(n93), .B(n91), .O(po02));
  invx g0051(.A(n92), .O(n91));
  orx  g0052(.A(n94), .B(n747), .O(n92));
  andx g0053(.A(n747), .B(n94), .O(n93));
  andx g0054(.A(n96), .B(n95), .O(n94));
  orx  g0055(.A(n98), .B(n753), .O(n95));
  invx g0056(.A(n97), .O(n96));
  andx g0057(.A(n753), .B(n98), .O(n97));
  invx g0058(.A(n752), .O(n98));
  orx  g0059(.A(n101), .B(n100), .O(po01));
  andx g0060(.A(n103), .B(n104), .O(n100));
  invx g0061(.A(n102), .O(n101));
  orx  g0062(.A(n104), .B(n103), .O(n102));
  andx g0063(.A(pi00), .B(pi03), .O(n103));
  orx  g0064(.A(n105), .B(n40), .O(n104));
  invx g0065(.A(pi01), .O(n105));
  orx  g0066(.A(n121), .B(n107), .O(po19));
  orx  g0067(.A(n109), .B(n108), .O(n107));
  andx g0068(.A(n114), .B(n116), .O(n108));
  invx g0069(.A(n113), .O(n109));
  orx  g0070(.A(n115), .B(n111), .O(po18));
  andx g0071(.A(n112), .B(n117), .O(n111));
  andx g0072(.A(n114), .B(n113), .O(n112));
  orx  g0073(.A(n120), .B(n128), .O(n113));
  invx g0074(.A(n119), .O(n114));
  andx g0075(.A(n119), .B(n116), .O(n115));
  invx g0076(.A(n117), .O(n116));
  andx g0077(.A(n118), .B(n138), .O(n117));
  orx  g0078(.A(n139), .B(n134), .O(n118));
  andx g0079(.A(n128), .B(n120), .O(n119));
  orx  g0080(.A(n122), .B(n121), .O(n120));
  andx g0081(.A(pi02), .B(n125), .O(n121));
  andx g0082(.A(n124), .B(n123), .O(n122));
  orx  g0083(.A(n501), .B(n840), .O(n123));
  invx g0084(.A(n125), .O(n124));
  orx  g0085(.A(n126), .B(n151), .O(n125));
  andx g0086(.A(n127), .B(pi04), .O(n126));
  andx g0087(.A(pi06), .B(n149), .O(n127));
  orx  g0088(.A(n144), .B(n129), .O(n128));
  invx g0089(.A(n157), .O(n129));
  andx g0090(.A(n132), .B(n131), .O(po17));
  orx  g0091(.A(n134), .B(n136), .O(n131));
  invx g0092(.A(n133), .O(n132));
  andx g0093(.A(n136), .B(n134), .O(n133));
  andx g0094(.A(n135), .B(n165), .O(n134));
  orx  g0095(.A(n171), .B(n163), .O(n135));
  orx  g0096(.A(n139), .B(n137), .O(n136));
  invx g0097(.A(n138), .O(n137));
  orx  g0098(.A(n140), .B(n175), .O(n138));
  andx g0099(.A(n175), .B(n140), .O(n139));
  andx g0100(.A(n143), .B(n141), .O(n140));
  invx g0101(.A(n142), .O(n141));
  andx g0102(.A(n144), .B(n157), .O(n142));
  orx  g0103(.A(n157), .B(n144), .O(n143));
  orx  g0104(.A(n147), .B(n145), .O(n144));
  invx g0105(.A(n146), .O(n145));
  orx  g0106(.A(n148), .B(n156), .O(n146));
  andx g0107(.A(n156), .B(n148), .O(n147));
  andx g0108(.A(n150), .B(n149), .O(n148));
  orx  g0109(.A(n152), .B(n155), .O(n149));
  invx g0110(.A(n151), .O(n150));
  andx g0111(.A(n155), .B(n152), .O(n151));
  orx  g0112(.A(n153), .B(n189), .O(n152));
  andx g0113(.A(n154), .B(pi04), .O(n153));
  andx g0114(.A(pi19), .B(n187), .O(n154));
  andx g0115(.A(pi07), .B(pi02), .O(n155));
  andx g0116(.A(pi06), .B(pi04), .O(n156));
  orx  g0117(.A(n158), .B(n196), .O(n157));
  andx g0118(.A(n182), .B(n159), .O(n158));
  orx  g0119(.A(n160), .B(n200), .O(n159));
  andx g0120(.A(pi02), .B(pi18), .O(n160));
  orx  g0121(.A(n167), .B(n162), .O(po16));
  andx g0122(.A(n164), .B(n163), .O(n162));
  invx g0123(.A(n168), .O(n163));
  andx g0124(.A(n172), .B(n165), .O(n164));
  invx g0125(.A(n166), .O(n165));
  andx g0126(.A(n173), .B(n206), .O(n166));
  andx g0127(.A(n171), .B(n168), .O(n167));
  orx  g0128(.A(n170), .B(n169), .O(n168));
  andx g0129(.A(n213), .B(n209), .O(n169));
  andx g0130(.A(n280), .B(n214), .O(n170));
  invx g0131(.A(n172), .O(n171));
  orx  g0132(.A(n206), .B(n173), .O(n172));
  andx g0133(.A(n175), .B(n174), .O(n173));
  orx  g0134(.A(n204), .B(n177), .O(n174));
  invx g0135(.A(n176), .O(n175));
  andx g0136(.A(n204), .B(n177), .O(n176));
  andx g0137(.A(n180), .B(n178), .O(n177));
  invx g0138(.A(n179), .O(n178));
  andx g0139(.A(n181), .B(n195), .O(n179));
  orx  g0140(.A(n195), .B(n181), .O(n180));
  invx g0141(.A(n182), .O(n181));
  andx g0142(.A(n184), .B(n183), .O(n182));
  orx  g0143(.A(n186), .B(n194), .O(n183));
  invx g0144(.A(n185), .O(n184));
  andx g0145(.A(n194), .B(n186), .O(n185));
  andx g0146(.A(n188), .B(n187), .O(n186));
  orx  g0147(.A(n190), .B(n193), .O(n187));
  invx g0148(.A(n189), .O(n188));
  andx g0149(.A(n193), .B(n190), .O(n189));
  orx  g0150(.A(n191), .B(n237), .O(n190));
  andx g0151(.A(n192), .B(pi04), .O(n191));
  andx g0152(.A(pi16), .B(n235), .O(n192));
  andx g0153(.A(pi06), .B(pi07), .O(n193));
  andx g0154(.A(pi19), .B(pi04), .O(n194));
  orx  g0155(.A(n197), .B(n196), .O(n195));
  andx g0156(.A(n200), .B(pi02), .O(n196));
  andx g0157(.A(n199), .B(n198), .O(n197));
  orx  g0158(.A(n992), .B(n501), .O(n198));
  invx g0159(.A(n200), .O(n199));
  orx  g0160(.A(n201), .B(n244), .O(n200));
  andx g0161(.A(n228), .B(n202), .O(n201));
  orx  g0162(.A(n203), .B(n248), .O(n202));
  andx g0163(.A(pi06), .B(pi18), .O(n203));
  orx  g0164(.A(n205), .B(n256), .O(n204));
  andx g0165(.A(n225), .B(n253), .O(n205));
  andx g0166(.A(n259), .B(n219), .O(n206));
  andx g0167(.A(n210), .B(n208), .O(po15));
  orx  g0168(.A(n212), .B(n209), .O(n208));
  invx g0169(.A(n263), .O(n209));
  orx  g0170(.A(n263), .B(n211), .O(n210));
  invx g0171(.A(n212), .O(n211));
  andx g0172(.A(n215), .B(n213), .O(n212));
  orx  g0173(.A(n280), .B(n214), .O(n213));
  invx g0174(.A(n216), .O(n214));
  orx  g0175(.A(n279), .B(n216), .O(n215));
  andx g0176(.A(n220), .B(n217), .O(n216));
  orx  g0177(.A(n219), .B(n218), .O(n217));
  invx g0178(.A(n259), .O(n218));
  invx g0179(.A(n221), .O(n219));
  orx  g0180(.A(n259), .B(n221), .O(n220));
  orx  g0181(.A(n224), .B(n222), .O(n221));
  invx g0182(.A(n223), .O(n222));
  orx  g0183(.A(n225), .B(n252), .O(n223));
  andx g0184(.A(n252), .B(n225), .O(n224));
  andx g0185(.A(n229), .B(n226), .O(n225));
  orx  g0186(.A(n228), .B(n227), .O(n226));
  invx g0187(.A(n243), .O(n227));
  invx g0188(.A(n230), .O(n228));
  orx  g0189(.A(n243), .B(n230), .O(n229));
  orx  g0190(.A(n233), .B(n231), .O(n230));
  invx g0191(.A(n232), .O(n231));
  orx  g0192(.A(n234), .B(n242), .O(n232));
  andx g0193(.A(n242), .B(n234), .O(n233));
  andx g0194(.A(n236), .B(n235), .O(n234));
  orx  g0195(.A(n238), .B(n241), .O(n235));
  invx g0196(.A(n237), .O(n236));
  andx g0197(.A(n241), .B(n238), .O(n237));
  orx  g0198(.A(n239), .B(n301), .O(n238));
  andx g0199(.A(n240), .B(pi04), .O(n239));
  andx g0200(.A(pi14), .B(n299), .O(n240));
  andx g0201(.A(pi19), .B(pi07), .O(n241));
  andx g0202(.A(pi16), .B(pi04), .O(n242));
  orx  g0203(.A(n245), .B(n244), .O(n243));
  andx g0204(.A(n248), .B(pi06), .O(n244));
  andx g0205(.A(n247), .B(n246), .O(n245));
  orx  g0206(.A(n992), .B(n895), .O(n246));
  invx g0207(.A(n248), .O(n247));
  orx  g0208(.A(n249), .B(n308), .O(n248));
  andx g0209(.A(n292), .B(n250), .O(n249));
  orx  g0210(.A(n251), .B(n312), .O(n250));
  andx g0211(.A(pi18), .B(pi19), .O(n251));
  andx g0212(.A(n255), .B(n253), .O(n252));
  orx  g0213(.A(n254), .B(n257), .O(n253));
  andx g0214(.A(pi02), .B(pi17), .O(n254));
  invx g0215(.A(n256), .O(n255));
  andx g0216(.A(n257), .B(pi02), .O(n256));
  orx  g0217(.A(n258), .B(n320), .O(n257));
  andx g0218(.A(n289), .B(n317), .O(n258));
  orx  g0219(.A(n260), .B(n325), .O(n259));
  andx g0220(.A(n285), .B(n261), .O(n260));
  orx  g0221(.A(n262), .B(n329), .O(n261));
  andx g0222(.A(pi02), .B(pi15), .O(n262));
  andx g0223(.A(n267), .B(n272), .O(n263));
  andx g0224(.A(n272), .B(n265), .O(po14));
  orx  g0225(.A(n266), .B(n274), .O(n265));
  andx g0226(.A(n270), .B(n267), .O(n266));
  orx  g0227(.A(n350), .B(n268), .O(n267));
  orx  g0228(.A(n347), .B(n269), .O(n268));
  invx g0229(.A(n277), .O(n269));
  orx  g0230(.A(n271), .B(n277), .O(n270));
  andx g0231(.A(n348), .B(n411), .O(n271));
  invx g0232(.A(n273), .O(n272));
  andx g0233(.A(n277), .B(n274), .O(n273));
  orx  g0234(.A(n275), .B(n342), .O(n274));
  invx g0235(.A(n276), .O(n275));
  orx  g0236(.A(n344), .B(n339), .O(n276));
  andx g0237(.A(n279), .B(n278), .O(n277));
  orx  g0238(.A(n333), .B(n281), .O(n278));
  invx g0239(.A(n280), .O(n279));
  andx g0240(.A(n333), .B(n281), .O(n280));
  andx g0241(.A(n283), .B(n282), .O(n281));
  orx  g0242(.A(n285), .B(n323), .O(n282));
  invx g0243(.A(n284), .O(n283));
  andx g0244(.A(n323), .B(n285), .O(n284));
  andx g0245(.A(n287), .B(n286), .O(n285));
  orx  g0246(.A(n289), .B(n316), .O(n286));
  invx g0247(.A(n288), .O(n287));
  andx g0248(.A(n316), .B(n289), .O(n288));
  andx g0249(.A(n293), .B(n290), .O(n289));
  orx  g0250(.A(n292), .B(n291), .O(n290));
  invx g0251(.A(n307), .O(n291));
  invx g0252(.A(n294), .O(n292));
  orx  g0253(.A(n307), .B(n294), .O(n293));
  orx  g0254(.A(n297), .B(n295), .O(n294));
  invx g0255(.A(n296), .O(n295));
  orx  g0256(.A(n298), .B(n306), .O(n296));
  andx g0257(.A(n306), .B(n298), .O(n297));
  andx g0258(.A(n300), .B(n299), .O(n298));
  orx  g0259(.A(n302), .B(n305), .O(n299));
  invx g0260(.A(n301), .O(n300));
  andx g0261(.A(n305), .B(n302), .O(n301));
  orx  g0262(.A(n303), .B(n375), .O(n302));
  andx g0263(.A(n304), .B(pi04), .O(n303));
  andx g0264(.A(pi13), .B(n373), .O(n304));
  andx g0265(.A(pi16), .B(pi07), .O(n305));
  andx g0266(.A(pi14), .B(pi04), .O(n306));
  orx  g0267(.A(n309), .B(n308), .O(n307));
  andx g0268(.A(n312), .B(pi19), .O(n308));
  andx g0269(.A(n311), .B(n310), .O(n309));
  orx  g0270(.A(n483), .B(n992), .O(n310));
  invx g0271(.A(n312), .O(n311));
  orx  g0272(.A(n313), .B(n382), .O(n312));
  andx g0273(.A(n366), .B(n314), .O(n313));
  orx  g0274(.A(n315), .B(n386), .O(n314));
  andx g0275(.A(pi18), .B(pi16), .O(n315));
  andx g0276(.A(n319), .B(n317), .O(n316));
  orx  g0277(.A(n318), .B(n321), .O(n317));
  andx g0278(.A(pi06), .B(pi17), .O(n318));
  invx g0279(.A(n320), .O(n319));
  andx g0280(.A(n321), .B(pi06), .O(n320));
  orx  g0281(.A(n322), .B(n392), .O(n321));
  andx g0282(.A(n363), .B(n389), .O(n322));
  invx g0283(.A(n324), .O(n323));
  orx  g0284(.A(n326), .B(n325), .O(n324));
  andx g0285(.A(n329), .B(pi02), .O(n325));
  andx g0286(.A(n328), .B(n327), .O(n326));
  orx  g0287(.A(n1160), .B(n501), .O(n327));
  invx g0288(.A(n329), .O(n328));
  orx  g0289(.A(n330), .B(n396), .O(n329));
  andx g0290(.A(n357), .B(n331), .O(n330));
  orx  g0291(.A(n332), .B(n400), .O(n331));
  andx g0292(.A(pi06), .B(pi15), .O(n332));
  orx  g0293(.A(n334), .B(n408), .O(n333));
  andx g0294(.A(n354), .B(n405), .O(n334));
  andx g0295(.A(n337), .B(n336), .O(po13));
  orx  g0296(.A(n339), .B(n341), .O(n336));
  invx g0297(.A(n338), .O(n337));
  andx g0298(.A(n341), .B(n339), .O(n338));
  andx g0299(.A(n340), .B(n420), .O(n339));
  orx  g0300(.A(n512), .B(n424), .O(n340));
  orx  g0301(.A(n344), .B(n342), .O(n341));
  invx g0302(.A(n343), .O(n342));
  orx  g0303(.A(n345), .B(n427), .O(n343));
  andx g0304(.A(n427), .B(n345), .O(n344));
  andx g0305(.A(n349), .B(n346), .O(n345));
  orx  g0306(.A(n348), .B(n347), .O(n346));
  invx g0307(.A(n411), .O(n347));
  invx g0308(.A(n350), .O(n348));
  orx  g0309(.A(n411), .B(n350), .O(n349));
  orx  g0310(.A(n353), .B(n351), .O(n350));
  invx g0311(.A(n352), .O(n351));
  orx  g0312(.A(n354), .B(n404), .O(n352));
  andx g0313(.A(n404), .B(n354), .O(n353));
  andx g0314(.A(n358), .B(n355), .O(n354));
  orx  g0315(.A(n357), .B(n356), .O(n355));
  invx g0316(.A(n395), .O(n356));
  invx g0317(.A(n359), .O(n357));
  orx  g0318(.A(n395), .B(n359), .O(n358));
  orx  g0319(.A(n362), .B(n360), .O(n359));
  invx g0320(.A(n361), .O(n360));
  orx  g0321(.A(n363), .B(n388), .O(n361));
  andx g0322(.A(n388), .B(n363), .O(n362));
  andx g0323(.A(n367), .B(n364), .O(n363));
  orx  g0324(.A(n366), .B(n365), .O(n364));
  invx g0325(.A(n381), .O(n365));
  invx g0326(.A(n368), .O(n366));
  orx  g0327(.A(n381), .B(n368), .O(n367));
  orx  g0328(.A(n371), .B(n369), .O(n368));
  invx g0329(.A(n370), .O(n369));
  orx  g0330(.A(n372), .B(n380), .O(n370));
  andx g0331(.A(n380), .B(n372), .O(n371));
  andx g0332(.A(n374), .B(n373), .O(n372));
  orx  g0333(.A(n376), .B(n379), .O(n373));
  invx g0334(.A(n375), .O(n374));
  andx g0335(.A(n379), .B(n376), .O(n375));
  orx  g0336(.A(n377), .B(n456), .O(n376));
  andx g0337(.A(n378), .B(pi04), .O(n377));
  andx g0338(.A(pi10), .B(n454), .O(n378));
  andx g0339(.A(pi14), .B(pi07), .O(n379));
  andx g0340(.A(pi13), .B(pi04), .O(n380));
  orx  g0341(.A(n383), .B(n382), .O(n381));
  andx g0342(.A(n386), .B(pi16), .O(n382));
  andx g0343(.A(n385), .B(n384), .O(n383));
  orx  g0344(.A(n1031), .B(n992), .O(n384));
  invx g0345(.A(n386), .O(n385));
  orx  g0346(.A(n387), .B(n465), .O(n386));
  andx g0347(.A(n449), .B(n466), .O(n387));
  andx g0348(.A(n391), .B(n389), .O(n388));
  orx  g0349(.A(n390), .B(n393), .O(n389));
  andx g0350(.A(pi19), .B(pi17), .O(n390));
  invx g0351(.A(n392), .O(n391));
  andx g0352(.A(n393), .B(pi19), .O(n392));
  orx  g0353(.A(n394), .B(n476), .O(n393));
  andx g0354(.A(n445), .B(n473), .O(n394));
  orx  g0355(.A(n397), .B(n396), .O(n395));
  andx g0356(.A(n400), .B(pi06), .O(n396));
  andx g0357(.A(n399), .B(n398), .O(n397));
  orx  g0358(.A(n895), .B(n1160), .O(n398));
  invx g0359(.A(n400), .O(n399));
  orx  g0360(.A(n401), .B(n480), .O(n400));
  andx g0361(.A(n439), .B(n402), .O(n401));
  orx  g0362(.A(n403), .B(n485), .O(n402));
  andx g0363(.A(pi19), .B(pi15), .O(n403));
  andx g0364(.A(n407), .B(n405), .O(n404));
  orx  g0365(.A(n406), .B(n409), .O(n405));
  andx g0366(.A(pi02), .B(pi12), .O(n406));
  invx g0367(.A(n408), .O(n407));
  andx g0368(.A(n409), .B(pi02), .O(n408));
  orx  g0369(.A(n410), .B(n493), .O(n409));
  andx g0370(.A(n436), .B(n490), .O(n410));
  orx  g0371(.A(n412), .B(n498), .O(n411));
  andx g0372(.A(n431), .B(n413), .O(n412));
  orx  g0373(.A(n414), .B(n503), .O(n413));
  andx g0374(.A(pi02), .B(pi11), .O(n414));
  orx  g0375(.A(n417), .B(n416), .O(po12));
  andx g0376(.A(n419), .B(n512), .O(n416));
  invx g0377(.A(n418), .O(n417));
  orx  g0378(.A(n512), .B(n419), .O(n418));
  andx g0379(.A(n422), .B(n420), .O(n419));
  orx  g0380(.A(n520), .B(n421), .O(n420));
  orx  g0381(.A(n608), .B(n424), .O(n421));
  invx g0382(.A(n423), .O(n422));
  andx g0383(.A(n510), .B(n424), .O(n423));
  orx  g0384(.A(n426), .B(n425), .O(n424));
  andx g0385(.A(n507), .B(n428), .O(n425));
  invx g0386(.A(n427), .O(n426));
  orx  g0387(.A(n507), .B(n428), .O(n427));
  orx  g0388(.A(n430), .B(n429), .O(n428));
  andx g0389(.A(n432), .B(n497), .O(n429));
  andx g0390(.A(n496), .B(n431), .O(n430));
  invx g0391(.A(n432), .O(n431));
  orx  g0392(.A(n435), .B(n433), .O(n432));
  invx g0393(.A(n434), .O(n433));
  orx  g0394(.A(n436), .B(n489), .O(n434));
  andx g0395(.A(n489), .B(n436), .O(n435));
  andx g0396(.A(n440), .B(n437), .O(n436));
  orx  g0397(.A(n439), .B(n438), .O(n437));
  invx g0398(.A(n479), .O(n438));
  invx g0399(.A(n441), .O(n439));
  orx  g0400(.A(n479), .B(n441), .O(n440));
  orx  g0401(.A(n444), .B(n442), .O(n441));
  invx g0402(.A(n443), .O(n442));
  orx  g0403(.A(n445), .B(n472), .O(n443));
  andx g0404(.A(n472), .B(n445), .O(n444));
  andx g0405(.A(n447), .B(n446), .O(n445));
  orx  g0406(.A(n449), .B(n463), .O(n446));
  invx g0407(.A(n448), .O(n447));
  andx g0408(.A(n463), .B(n449), .O(n448));
  andx g0409(.A(n451), .B(n450), .O(n449));
  orx  g0410(.A(n453), .B(n462), .O(n450));
  invx g0411(.A(n452), .O(n451));
  andx g0412(.A(n462), .B(n453), .O(n452));
  andx g0413(.A(n455), .B(n454), .O(n453));
  orx  g0414(.A(n457), .B(n461), .O(n454));
  invx g0415(.A(n456), .O(n455));
  andx g0416(.A(n461), .B(n457), .O(n456));
  orx  g0417(.A(n459), .B(n458), .O(n457));
  andx g0418(.A(n556), .B(n559), .O(n458));
  andx g0419(.A(n460), .B(n557), .O(n459));
  orx  g0420(.A(n559), .B(n556), .O(n460));
  andx g0421(.A(pi13), .B(pi07), .O(n461));
  andx g0422(.A(pi10), .B(pi04), .O(n462));
  andx g0423(.A(n466), .B(n464), .O(n463));
  invx g0424(.A(n465), .O(n464));
  andx g0425(.A(n468), .B(pi14), .O(n465));
  orx  g0426(.A(n468), .B(n467), .O(n466));
  andx g0427(.A(pi14), .B(pi18), .O(n467));
  orx  g0428(.A(n469), .B(n561), .O(n468));
  andx g0429(.A(n547), .B(n470), .O(n469));
  orx  g0430(.A(n471), .B(n565), .O(n470));
  andx g0431(.A(pi18), .B(pi13), .O(n471));
  andx g0432(.A(n475), .B(n473), .O(n472));
  orx  g0433(.A(n474), .B(n477), .O(n473));
  andx g0434(.A(pi17), .B(pi16), .O(n474));
  invx g0435(.A(n476), .O(n475));
  andx g0436(.A(n477), .B(pi16), .O(n476));
  orx  g0437(.A(n478), .B(n571), .O(n477));
  andx g0438(.A(n542), .B(n568), .O(n478));
  orx  g0439(.A(n481), .B(n480), .O(n479));
  andx g0440(.A(n485), .B(pi19), .O(n480));
  andx g0441(.A(n484), .B(n482), .O(n481));
  orx  g0442(.A(n1160), .B(n483), .O(n482));
  invx g0443(.A(pi19), .O(n483));
  invx g0444(.A(n485), .O(n484));
  orx  g0445(.A(n486), .B(n577), .O(n485));
  andx g0446(.A(n536), .B(n487), .O(n486));
  orx  g0447(.A(n488), .B(n581), .O(n487));
  andx g0448(.A(pi16), .B(pi15), .O(n488));
  andx g0449(.A(n492), .B(n490), .O(n489));
  orx  g0450(.A(n491), .B(n494), .O(n490));
  andx g0451(.A(pi06), .B(pi12), .O(n491));
  invx g0452(.A(n493), .O(n492));
  andx g0453(.A(n494), .B(pi06), .O(n493));
  orx  g0454(.A(n495), .B(n587), .O(n494));
  andx g0455(.A(n533), .B(n584), .O(n495));
  invx g0456(.A(n497), .O(n496));
  orx  g0457(.A(n499), .B(n498), .O(n497));
  andx g0458(.A(n503), .B(pi02), .O(n498));
  andx g0459(.A(n502), .B(n500), .O(n499));
  orx  g0460(.A(n1137), .B(n501), .O(n500));
  invx g0461(.A(pi02), .O(n501));
  invx g0462(.A(n503), .O(n502));
  orx  g0463(.A(n504), .B(n593), .O(n503));
  andx g0464(.A(n527), .B(n505), .O(n504));
  orx  g0465(.A(n506), .B(n597), .O(n505));
  andx g0466(.A(pi06), .B(pi11), .O(n506));
  andx g0467(.A(n508), .B(n602), .O(n507));
  invx g0468(.A(n509), .O(n508));
  andx g0469(.A(n524), .B(n600), .O(n509));
  orx  g0470(.A(n608), .B(n520), .O(n510));
  andx g0471(.A(n515), .B(n512), .O(po11));
  orx  g0472(.A(n616), .B(n513), .O(n512));
  invx g0473(.A(n514), .O(n513));
  andx g0474(.A(n715), .B(n516), .O(n514));
  orx  g0475(.A(n611), .B(n516), .O(n515));
  orx  g0476(.A(n518), .B(n517), .O(n516));
  andx g0477(.A(n520), .B(n609), .O(n517));
  andx g0478(.A(n608), .B(n519), .O(n518));
  invx g0479(.A(n520), .O(n519));
  orx  g0480(.A(n523), .B(n521), .O(n520));
  invx g0481(.A(n522), .O(n521));
  orx  g0482(.A(n524), .B(n599), .O(n522));
  andx g0483(.A(n599), .B(n524), .O(n523));
  andx g0484(.A(n528), .B(n525), .O(n524));
  orx  g0485(.A(n527), .B(n526), .O(n525));
  invx g0486(.A(n592), .O(n526));
  invx g0487(.A(n529), .O(n527));
  orx  g0488(.A(n592), .B(n529), .O(n528));
  orx  g0489(.A(n532), .B(n530), .O(n529));
  invx g0490(.A(n531), .O(n530));
  orx  g0491(.A(n533), .B(n583), .O(n531));
  andx g0492(.A(n583), .B(n533), .O(n532));
  andx g0493(.A(n537), .B(n534), .O(n533));
  orx  g0494(.A(n536), .B(n535), .O(n534));
  invx g0495(.A(n576), .O(n535));
  invx g0496(.A(n538), .O(n536));
  orx  g0497(.A(n576), .B(n538), .O(n537));
  orx  g0498(.A(n541), .B(n539), .O(n538));
  invx g0499(.A(n540), .O(n539));
  orx  g0500(.A(n542), .B(n567), .O(n540));
  andx g0501(.A(n567), .B(n542), .O(n541));
  andx g0502(.A(n545), .B(n543), .O(n542));
  orx  g0503(.A(n547), .B(n544), .O(n543));
  invx g0504(.A(n560), .O(n544));
  orx  g0505(.A(n560), .B(n546), .O(n545));
  invx g0506(.A(n547), .O(n546));
  andx g0507(.A(n550), .B(n548), .O(n547));
  invx g0508(.A(n549), .O(n548));
  andx g0509(.A(n551), .B(n557), .O(n549));
  orx  g0510(.A(n557), .B(n551), .O(n550));
  orx  g0511(.A(n554), .B(n552), .O(n551));
  andx g0512(.A(n559), .B(n553), .O(n552));
  invx g0513(.A(n556), .O(n553));
  andx g0514(.A(n556), .B(n555), .O(n554));
  invx g0515(.A(n559), .O(n555));
  andx g0516(.A(pi10), .B(pi07), .O(n556));
  orx  g0517(.A(n558), .B(n653), .O(n557));
  andx g0518(.A(n559), .B(n841), .O(n558));
  andx g0519(.A(pi08), .B(pi04), .O(n559));
  orx  g0520(.A(n562), .B(n561), .O(n560));
  andx g0521(.A(n565), .B(pi13), .O(n561));
  andx g0522(.A(n564), .B(n563), .O(n562));
  orx  g0523(.A(n1117), .B(n992), .O(n563));
  invx g0524(.A(n565), .O(n564));
  orx  g0525(.A(n566), .B(n660), .O(n565));
  andx g0526(.A(n645), .B(n658), .O(n566));
  andx g0527(.A(n570), .B(n568), .O(n567));
  orx  g0528(.A(n569), .B(n572), .O(n568));
  andx g0529(.A(pi17), .B(pi14), .O(n569));
  invx g0530(.A(n571), .O(n570));
  andx g0531(.A(n572), .B(pi14), .O(n571));
  orx  g0532(.A(n573), .B(n668), .O(n572));
  andx g0533(.A(n641), .B(n574), .O(n573));
  orx  g0534(.A(n575), .B(n672), .O(n574));
  andx g0535(.A(pi17), .B(pi13), .O(n575));
  orx  g0536(.A(n578), .B(n577), .O(n576));
  andx g0537(.A(n581), .B(pi16), .O(n577));
  andx g0538(.A(n580), .B(n579), .O(n578));
  orx  g0539(.A(n1160), .B(n1031), .O(n579));
  invx g0540(.A(n581), .O(n580));
  orx  g0541(.A(n582), .B(n678), .O(n581));
  andx g0542(.A(n637), .B(n676), .O(n582));
  andx g0543(.A(n586), .B(n584), .O(n583));
  orx  g0544(.A(n585), .B(n588), .O(n584));
  andx g0545(.A(pi19), .B(pi12), .O(n585));
  invx g0546(.A(n587), .O(n586));
  andx g0547(.A(n588), .B(pi19), .O(n587));
  orx  g0548(.A(n589), .B(n684), .O(n588));
  andx g0549(.A(n633), .B(n590), .O(n589));
  orx  g0550(.A(n591), .B(n688), .O(n590));
  andx g0551(.A(pi16), .B(pi12), .O(n591));
  orx  g0552(.A(n594), .B(n593), .O(n592));
  andx g0553(.A(n597), .B(pi06), .O(n593));
  andx g0554(.A(n596), .B(n595), .O(n594));
  orx  g0555(.A(n1137), .B(n895), .O(n595));
  invx g0556(.A(n597), .O(n596));
  orx  g0557(.A(n598), .B(n694), .O(n597));
  andx g0558(.A(n629), .B(n692), .O(n598));
  andx g0559(.A(n602), .B(n600), .O(n599));
  orx  g0560(.A(n601), .B(n604), .O(n600));
  andx g0561(.A(pi02), .B(pi09), .O(n601));
  invx g0562(.A(n603), .O(n602));
  andx g0563(.A(n604), .B(pi02), .O(n603));
  orx  g0564(.A(n605), .B(n700), .O(n604));
  andx g0565(.A(n625), .B(n606), .O(n605));
  orx  g0566(.A(n607), .B(n704), .O(n606));
  andx g0567(.A(pi06), .B(pi09), .O(n607));
  invx g0568(.A(n609), .O(n608));
  orx  g0569(.A(n610), .B(n710), .O(n609));
  andx g0570(.A(n621), .B(n707), .O(n610));
  andx g0571(.A(n617), .B(n715), .O(n611));
  orx  g0572(.A(n614), .B(n613), .O(po10));
  andx g0573(.A(n616), .B(n715), .O(n613));
  invx g0574(.A(n615), .O(n614));
  orx  g0575(.A(n715), .B(n616), .O(n615));
  invx g0576(.A(n617), .O(n616));
  andx g0577(.A(n619), .B(n618), .O(n617));
  orx  g0578(.A(n621), .B(n706), .O(n618));
  invx g0579(.A(n620), .O(n619));
  andx g0580(.A(n706), .B(n621), .O(n620));
  orx  g0581(.A(n623), .B(n622), .O(n621));
  andx g0582(.A(n625), .B(n699), .O(n622));
  invx g0583(.A(n624), .O(n623));
  orx  g0584(.A(n699), .B(n625), .O(n624));
  orx  g0585(.A(n627), .B(n626), .O(n625));
  andx g0586(.A(n629), .B(n690), .O(n626));
  invx g0587(.A(n628), .O(n627));
  orx  g0588(.A(n690), .B(n629), .O(n628));
  orx  g0589(.A(n631), .B(n630), .O(n629));
  andx g0590(.A(n633), .B(n683), .O(n630));
  invx g0591(.A(n632), .O(n631));
  orx  g0592(.A(n683), .B(n633), .O(n632));
  orx  g0593(.A(n635), .B(n634), .O(n633));
  andx g0594(.A(n637), .B(n674), .O(n634));
  invx g0595(.A(n636), .O(n635));
  orx  g0596(.A(n674), .B(n637), .O(n636));
  orx  g0597(.A(n639), .B(n638), .O(n637));
  andx g0598(.A(n641), .B(n667), .O(n638));
  invx g0599(.A(n640), .O(n639));
  orx  g0600(.A(n667), .B(n641), .O(n640));
  orx  g0601(.A(n643), .B(n642), .O(n641));
  andx g0602(.A(n645), .B(n656), .O(n642));
  invx g0603(.A(n644), .O(n643));
  orx  g0604(.A(n656), .B(n645), .O(n644));
  orx  g0605(.A(n647), .B(n646), .O(n645));
  andx g0606(.A(n649), .B(n655), .O(n646));
  invx g0607(.A(n648), .O(n647));
  orx  g0608(.A(n655), .B(n649), .O(n648));
  orx  g0609(.A(n652), .B(n650), .O(n649));
  andx g0610(.A(n651), .B(pi08), .O(n650));
  andx g0611(.A(pi07), .B(n654), .O(n651));
  andx g0612(.A(n653), .B(n848), .O(n652));
  invx g0613(.A(n654), .O(n653));
  orx  g0614(.A(n840), .B(n846), .O(n654));
  orx  g0615(.A(n40), .B(n840), .O(n655));
  orx  g0616(.A(n660), .B(n657), .O(n656));
  invx g0617(.A(n658), .O(n657));
  orx  g0618(.A(n659), .B(n661), .O(n658));
  andx g0619(.A(pi18), .B(pi10), .O(n659));
  andx g0620(.A(n661), .B(pi10), .O(n660));
  orx  g0621(.A(n664), .B(n662), .O(n661));
  andx g0622(.A(n663), .B(pi18), .O(n662));
  andx g0623(.A(pi08), .B(n835), .O(n663));
  andx g0624(.A(n665), .B(n1000), .O(n664));
  andx g0625(.A(n1001), .B(n666), .O(n665));
  orx  g0626(.A(pi08), .B(n835), .O(n666));
  orx  g0627(.A(n669), .B(n668), .O(n667));
  andx g0628(.A(n672), .B(pi13), .O(n668));
  andx g0629(.A(n671), .B(n670), .O(n669));
  orx  g0630(.A(n1117), .B(n1103), .O(n670));
  invx g0631(.A(n672), .O(n671));
  orx  g0632(.A(n673), .B(n854), .O(n672));
  andx g0633(.A(n831), .B(n852), .O(n673));
  orx  g0634(.A(n678), .B(n675), .O(n674));
  invx g0635(.A(n676), .O(n675));
  orx  g0636(.A(n677), .B(n679), .O(n676));
  andx g0637(.A(pi15), .B(pi14), .O(n677));
  andx g0638(.A(n679), .B(pi14), .O(n678));
  orx  g0639(.A(n680), .B(n860), .O(n679));
  andx g0640(.A(n827), .B(n681), .O(n680));
  orx  g0641(.A(n682), .B(n864), .O(n681));
  andx g0642(.A(pi15), .B(pi13), .O(n682));
  orx  g0643(.A(n685), .B(n684), .O(n683));
  andx g0644(.A(n688), .B(pi16), .O(n684));
  andx g0645(.A(n687), .B(n686), .O(n685));
  orx  g0646(.A(n1149), .B(n1031), .O(n686));
  invx g0647(.A(n688), .O(n687));
  orx  g0648(.A(n689), .B(n870), .O(n688));
  andx g0649(.A(n823), .B(n868), .O(n689));
  orx  g0650(.A(n694), .B(n691), .O(n690));
  invx g0651(.A(n692), .O(n691));
  orx  g0652(.A(n693), .B(n695), .O(n692));
  andx g0653(.A(pi19), .B(pi11), .O(n693));
  andx g0654(.A(n695), .B(pi19), .O(n694));
  orx  g0655(.A(n696), .B(n876), .O(n695));
  andx g0656(.A(n819), .B(n697), .O(n696));
  orx  g0657(.A(n698), .B(n880), .O(n697));
  andx g0658(.A(pi16), .B(pi11), .O(n698));
  orx  g0659(.A(n701), .B(n700), .O(n699));
  andx g0660(.A(n704), .B(pi06), .O(n700));
  andx g0661(.A(n703), .B(n702), .O(n701));
  orx  g0662(.A(n1059), .B(n895), .O(n702));
  invx g0663(.A(n704), .O(n703));
  orx  g0664(.A(n705), .B(n886), .O(n704));
  andx g0665(.A(n815), .B(n884), .O(n705));
  andx g0666(.A(n709), .B(n707), .O(n706));
  orx  g0667(.A(n708), .B(n711), .O(n707));
  andx g0668(.A(pi02), .B(pi03), .O(n708));
  invx g0669(.A(n710), .O(n709));
  andx g0670(.A(n711), .B(pi02), .O(n710));
  orx  g0671(.A(n712), .B(n892), .O(n711));
  andx g0672(.A(n811), .B(n713), .O(n712));
  orx  g0673(.A(n714), .B(n897), .O(n713));
  andx g0674(.A(pi06), .B(pi03), .O(n714));
  orx  g0675(.A(n717), .B(n716), .O(n715));
  andx g0676(.A(n719), .B(pi02), .O(n716));
  andx g0677(.A(n807), .B(n718), .O(n717));
  orx  g0678(.A(n806), .B(n719), .O(n718));
  orx  g0679(.A(n721), .B(n720), .O(n719));
  andx g0680(.A(n723), .B(pi06), .O(n720));
  andx g0681(.A(n799), .B(n722), .O(n721));
  orx  g0682(.A(n798), .B(n723), .O(n722));
  orx  g0683(.A(n725), .B(n724), .O(n723));
  andx g0684(.A(n727), .B(pi19), .O(n724));
  andx g0685(.A(n790), .B(n726), .O(n725));
  orx  g0686(.A(n789), .B(n727), .O(n726));
  orx  g0687(.A(n729), .B(n728), .O(n727));
  andx g0688(.A(n731), .B(pi16), .O(n728));
  andx g0689(.A(n782), .B(n730), .O(n729));
  orx  g0690(.A(n781), .B(n731), .O(n730));
  orx  g0691(.A(n733), .B(n732), .O(n731));
  andx g0692(.A(n735), .B(pi14), .O(n732));
  andx g0693(.A(n773), .B(n734), .O(n733));
  orx  g0694(.A(n772), .B(n735), .O(n734));
  orx  g0695(.A(n737), .B(n736), .O(n735));
  andx g0696(.A(n739), .B(pi13), .O(n736));
  andx g0697(.A(n765), .B(n738), .O(n737));
  orx  g0698(.A(n764), .B(n739), .O(n738));
  orx  g0699(.A(n741), .B(n740), .O(n739));
  andx g0700(.A(n743), .B(pi10), .O(n740));
  andx g0701(.A(n756), .B(n742), .O(n741));
  orx  g0702(.A(n755), .B(n743), .O(n742));
  orx  g0703(.A(n745), .B(n744), .O(n743));
  andx g0704(.A(n752), .B(n747), .O(n744));
  andx g0705(.A(n753), .B(n746), .O(n745));
  orx  g0706(.A(n752), .B(n747), .O(n746));
  orx  g0707(.A(n750), .B(n748), .O(n747));
  invx g0708(.A(n749), .O(n748));
  orx  g0709(.A(n751), .B(n754), .O(n749));
  andx g0710(.A(n754), .B(n751), .O(n750));
  orx  g0711(.A(n1151), .B(n1059), .O(n751));
  andx g0712(.A(pi01), .B(pi08), .O(n752));
  andx g0713(.A(n754), .B(po00), .O(n753));
  andx g0714(.A(pi05), .B(pi03), .O(n754));
  andx g0715(.A(pi10), .B(pi01), .O(n755));
  orx  g0716(.A(n759), .B(n757), .O(n756));
  invx g0717(.A(n758), .O(n757));
  orx  g0718(.A(n760), .B(n921), .O(n758));
  andx g0719(.A(n921), .B(n760), .O(n759));
  andx g0720(.A(n762), .B(n761), .O(n760));
  orx  g0721(.A(n929), .B(n927), .O(n761));
  orx  g0722(.A(n763), .B(n928), .O(n762));
  invx g0723(.A(n927), .O(n763));
  andx g0724(.A(pi13), .B(pi01), .O(n764));
  invx g0725(.A(n766), .O(n765));
  orx  g0726(.A(n768), .B(n767), .O(n766));
  andx g0727(.A(n770), .B(n933), .O(n767));
  invx g0728(.A(n769), .O(n768));
  orx  g0729(.A(n933), .B(n770), .O(n769));
  andx g0730(.A(n916), .B(n771), .O(n770));
  invx g0731(.A(n914), .O(n771));
  andx g0732(.A(pi14), .B(pi01), .O(n772));
  orx  g0733(.A(n775), .B(n774), .O(n773));
  andx g0734(.A(n942), .B(n777), .O(n774));
  invx g0735(.A(n776), .O(n775));
  orx  g0736(.A(n777), .B(n942), .O(n776));
  orx  g0737(.A(n778), .B(n910), .O(n777));
  andx g0738(.A(n780), .B(n779), .O(n778));
  orx  g0739(.A(n931), .B(n1117), .O(n779));
  invx g0740(.A(n913), .O(n780));
  andx g0741(.A(pi16), .B(pi01), .O(n781));
  invx g0742(.A(n783), .O(n782));
  orx  g0743(.A(n785), .B(n784), .O(n783));
  andx g0744(.A(n787), .B(n949), .O(n784));
  invx g0745(.A(n786), .O(n785));
  orx  g0746(.A(n949), .B(n787), .O(n786));
  andx g0747(.A(n908), .B(n788), .O(n787));
  invx g0748(.A(n906), .O(n788));
  andx g0749(.A(pi19), .B(pi01), .O(n789));
  orx  g0750(.A(n792), .B(n791), .O(n790));
  andx g0751(.A(n958), .B(n794), .O(n791));
  invx g0752(.A(n793), .O(n792));
  orx  g0753(.A(n794), .B(n958), .O(n793));
  orx  g0754(.A(n795), .B(n902), .O(n794));
  andx g0755(.A(n797), .B(n796), .O(n795));
  orx  g0756(.A(n931), .B(n1031), .O(n796));
  invx g0757(.A(n905), .O(n797));
  andx g0758(.A(pi06), .B(pi01), .O(n798));
  invx g0759(.A(n800), .O(n799));
  orx  g0760(.A(n802), .B(n801), .O(n800));
  andx g0761(.A(n804), .B(n965), .O(n801));
  invx g0762(.A(n803), .O(n802));
  orx  g0763(.A(n965), .B(n804), .O(n803));
  andx g0764(.A(n900), .B(n805), .O(n804));
  invx g0765(.A(n898), .O(n805));
  andx g0766(.A(pi02), .B(pi01), .O(n806));
  orx  g0767(.A(n809), .B(n808), .O(n807));
  andx g0768(.A(n811), .B(n891), .O(n808));
  invx g0769(.A(n810), .O(n809));
  orx  g0770(.A(n891), .B(n811), .O(n810));
  orx  g0771(.A(n813), .B(n812), .O(n811));
  andx g0772(.A(n815), .B(n882), .O(n812));
  invx g0773(.A(n814), .O(n813));
  orx  g0774(.A(n882), .B(n815), .O(n814));
  orx  g0775(.A(n817), .B(n816), .O(n815));
  andx g0776(.A(n819), .B(n875), .O(n816));
  invx g0777(.A(n818), .O(n817));
  orx  g0778(.A(n875), .B(n819), .O(n818));
  orx  g0779(.A(n821), .B(n820), .O(n819));
  andx g0780(.A(n823), .B(n866), .O(n820));
  invx g0781(.A(n822), .O(n821));
  orx  g0782(.A(n866), .B(n823), .O(n822));
  orx  g0783(.A(n825), .B(n824), .O(n823));
  andx g0784(.A(n827), .B(n859), .O(n824));
  invx g0785(.A(n826), .O(n825));
  orx  g0786(.A(n859), .B(n827), .O(n826));
  orx  g0787(.A(n829), .B(n828), .O(n827));
  andx g0788(.A(n831), .B(n850), .O(n828));
  invx g0789(.A(n830), .O(n829));
  orx  g0790(.A(n850), .B(n831), .O(n830));
  orx  g0791(.A(n833), .B(n832), .O(n831));
  andx g0792(.A(n835), .B(n842), .O(n832));
  invx g0793(.A(n834), .O(n833));
  orx  g0794(.A(n842), .B(n835), .O(n834));
  orx  g0795(.A(n838), .B(n836), .O(n835));
  invx g0796(.A(n837), .O(n836));
  orx  g0797(.A(n839), .B(n841), .O(n837));
  andx g0798(.A(n841), .B(n839), .O(n838));
  orx  g0799(.A(n1151), .B(n840), .O(n839));
  invx g0800(.A(pi04), .O(n840));
  andx g0801(.A(pi05), .B(pi07), .O(n841));
  invx g0802(.A(n843), .O(n842));
  orx  g0803(.A(n847), .B(n844), .O(n843));
  andx g0804(.A(n845), .B(pi08), .O(n844));
  andx g0805(.A(pi18), .B(n846), .O(n845));
  orx  g0806(.A(n1161), .B(n997), .O(n846));
  andx g0807(.A(n849), .B(n848), .O(n847));
  invx g0808(.A(pi08), .O(n848));
  andx g0809(.A(n1000), .B(n1001), .O(n849));
  orx  g0810(.A(n854), .B(n851), .O(n850));
  invx g0811(.A(n852), .O(n851));
  orx  g0812(.A(n853), .B(n855), .O(n852));
  andx g0813(.A(pi17), .B(pi10), .O(n853));
  andx g0814(.A(n855), .B(pi10), .O(n854));
  orx  g0815(.A(n857), .B(n856), .O(n855));
  andx g0816(.A(n994), .B(n995), .O(n856));
  andx g0817(.A(n989), .B(n858), .O(n857));
  orx  g0818(.A(n994), .B(n995), .O(n858));
  orx  g0819(.A(n861), .B(n860), .O(n859));
  andx g0820(.A(n864), .B(pi13), .O(n860));
  andx g0821(.A(n863), .B(n862), .O(n861));
  orx  g0822(.A(n1117), .B(n1160), .O(n862));
  invx g0823(.A(n864), .O(n863));
  orx  g0824(.A(n865), .B(n1006), .O(n864));
  andx g0825(.A(n982), .B(n1004), .O(n865));
  orx  g0826(.A(n870), .B(n867), .O(n866));
  invx g0827(.A(n868), .O(n867));
  orx  g0828(.A(n869), .B(n871), .O(n868));
  andx g0829(.A(pi14), .B(pi12), .O(n869));
  andx g0830(.A(n871), .B(pi14), .O(n870));
  orx  g0831(.A(n872), .B(n1012), .O(n871));
  andx g0832(.A(n978), .B(n873), .O(n872));
  orx  g0833(.A(n874), .B(n1016), .O(n873));
  andx g0834(.A(pi12), .B(pi13), .O(n874));
  orx  g0835(.A(n877), .B(n876), .O(n875));
  andx g0836(.A(n880), .B(pi16), .O(n876));
  andx g0837(.A(n879), .B(n878), .O(n877));
  orx  g0838(.A(n1137), .B(n1031), .O(n878));
  invx g0839(.A(n880), .O(n879));
  orx  g0840(.A(n881), .B(n1022), .O(n880));
  andx g0841(.A(n974), .B(n1020), .O(n881));
  orx  g0842(.A(n886), .B(n883), .O(n882));
  invx g0843(.A(n884), .O(n883));
  orx  g0844(.A(n885), .B(n887), .O(n884));
  andx g0845(.A(pi19), .B(pi09), .O(n885));
  andx g0846(.A(n887), .B(pi19), .O(n886));
  orx  g0847(.A(n888), .B(n1028), .O(n887));
  andx g0848(.A(n970), .B(n889), .O(n888));
  orx  g0849(.A(n890), .B(n1033), .O(n889));
  andx g0850(.A(pi16), .B(pi09), .O(n890));
  orx  g0851(.A(n893), .B(n892), .O(n891));
  andx g0852(.A(n897), .B(pi06), .O(n892));
  andx g0853(.A(n896), .B(n894), .O(n893));
  orx  g0854(.A(n931), .B(n895), .O(n894));
  invx g0855(.A(pi06), .O(n895));
  invx g0856(.A(n897), .O(n896));
  orx  g0857(.A(n899), .B(n898), .O(n897));
  andx g0858(.A(n901), .B(pi19), .O(n898));
  andx g0859(.A(n965), .B(n900), .O(n899));
  orx  g0860(.A(n964), .B(n901), .O(n900));
  orx  g0861(.A(n903), .B(n902), .O(n901));
  andx g0862(.A(n905), .B(pi16), .O(n902));
  andx g0863(.A(n958), .B(n904), .O(n903));
  orx  g0864(.A(n957), .B(n905), .O(n904));
  orx  g0865(.A(n907), .B(n906), .O(n905));
  andx g0866(.A(n909), .B(pi14), .O(n906));
  andx g0867(.A(n949), .B(n908), .O(n907));
  orx  g0868(.A(n948), .B(n909), .O(n908));
  orx  g0869(.A(n911), .B(n910), .O(n909));
  andx g0870(.A(n913), .B(pi13), .O(n910));
  andx g0871(.A(n942), .B(n912), .O(n911));
  orx  g0872(.A(n941), .B(n913), .O(n912));
  orx  g0873(.A(n915), .B(n914), .O(n913));
  andx g0874(.A(n917), .B(pi10), .O(n914));
  andx g0875(.A(n933), .B(n916), .O(n915));
  orx  g0876(.A(n932), .B(n917), .O(n916));
  orx  g0877(.A(n919), .B(n918), .O(n917));
  andx g0878(.A(n927), .B(n921), .O(n918));
  andx g0879(.A(n928), .B(n920), .O(n919));
  orx  g0880(.A(n927), .B(n921), .O(n920));
  orx  g0881(.A(n923), .B(n922), .O(n921));
  andx g0882(.A(n925), .B(n926), .O(n922));
  invx g0883(.A(n924), .O(n923));
  orx  g0884(.A(n926), .B(n925), .O(n924));
  andx g0885(.A(pi00), .B(pi11), .O(n925));
  orx  g0886(.A(n1161), .B(n1059), .O(n926));
  andx g0887(.A(pi03), .B(pi08), .O(n927));
  invx g0888(.A(n929), .O(n928));
  orx  g0889(.A(n41), .B(n930), .O(n929));
  orx  g0890(.A(n931), .B(n1059), .O(n930));
  invx g0891(.A(pi03), .O(n931));
  andx g0892(.A(pi10), .B(pi03), .O(n932));
  orx  g0893(.A(n936), .B(n934), .O(n933));
  invx g0894(.A(n935), .O(n934));
  orx  g0895(.A(n937), .B(n1049), .O(n935));
  andx g0896(.A(n1049), .B(n937), .O(n936));
  andx g0897(.A(n939), .B(n938), .O(n937));
  orx  g0898(.A(n1057), .B(n1055), .O(n938));
  orx  g0899(.A(n940), .B(n1056), .O(n939));
  invx g0900(.A(n1055), .O(n940));
  andx g0901(.A(pi13), .B(pi03), .O(n941));
  orx  g0902(.A(n944), .B(n943), .O(n942));
  andx g0903(.A(n1061), .B(n946), .O(n943));
  invx g0904(.A(n945), .O(n944));
  orx  g0905(.A(n946), .B(n1061), .O(n945));
  orx  g0906(.A(n1042), .B(n947), .O(n946));
  invx g0907(.A(n1044), .O(n947));
  andx g0908(.A(pi14), .B(pi03), .O(n948));
  orx  g0909(.A(n951), .B(n950), .O(n949));
  andx g0910(.A(n1070), .B(n953), .O(n950));
  invx g0911(.A(n952), .O(n951));
  orx  g0912(.A(n953), .B(n1070), .O(n952));
  orx  g0913(.A(n954), .B(n1038), .O(n953));
  andx g0914(.A(n956), .B(n955), .O(n954));
  orx  g0915(.A(n1059), .B(n1117), .O(n955));
  invx g0916(.A(n1041), .O(n956));
  andx g0917(.A(pi16), .B(pi03), .O(n957));
  orx  g0918(.A(n960), .B(n959), .O(n958));
  andx g0919(.A(n1077), .B(n962), .O(n959));
  invx g0920(.A(n961), .O(n960));
  orx  g0921(.A(n962), .B(n1077), .O(n961));
  orx  g0922(.A(n1034), .B(n963), .O(n962));
  invx g0923(.A(n1036), .O(n963));
  andx g0924(.A(pi19), .B(pi03), .O(n964));
  invx g0925(.A(n966), .O(n965));
  andx g0926(.A(n969), .B(n967), .O(n966));
  invx g0927(.A(n968), .O(n967));
  andx g0928(.A(n970), .B(n1027), .O(n968));
  orx  g0929(.A(n1027), .B(n970), .O(n969));
  orx  g0930(.A(n972), .B(n971), .O(n970));
  andx g0931(.A(n974), .B(n1018), .O(n971));
  invx g0932(.A(n973), .O(n972));
  orx  g0933(.A(n1018), .B(n974), .O(n973));
  orx  g0934(.A(n976), .B(n975), .O(n974));
  andx g0935(.A(n978), .B(n1011), .O(n975));
  invx g0936(.A(n977), .O(n976));
  orx  g0937(.A(n1011), .B(n978), .O(n977));
  orx  g0938(.A(n980), .B(n979), .O(n978));
  andx g0939(.A(n982), .B(n1002), .O(n979));
  invx g0940(.A(n981), .O(n980));
  orx  g0941(.A(n1002), .B(n982), .O(n981));
  orx  g0942(.A(n985), .B(n983), .O(n982));
  invx g0943(.A(n984), .O(n983));
  orx  g0944(.A(n986), .B(n995), .O(n984));
  andx g0945(.A(n995), .B(n986), .O(n985));
  andx g0946(.A(n988), .B(n987), .O(n986));
  orx  g0947(.A(n990), .B(n994), .O(n987));
  orx  g0948(.A(n993), .B(n989), .O(n988));
  invx g0949(.A(n990), .O(n989));
  orx  g0950(.A(n992), .B(n991), .O(n990));
  orx  g0951(.A(n41), .B(n1103), .O(n991));
  invx g0952(.A(pi18), .O(n992));
  invx g0953(.A(n994), .O(n993));
  andx g0954(.A(pi08), .B(pi17), .O(n994));
  orx  g0955(.A(n998), .B(n996), .O(n995));
  andx g0956(.A(n1000), .B(n997), .O(n996));
  invx g0957(.A(n1001), .O(n997));
  andx g0958(.A(n1001), .B(n999), .O(n998));
  invx g0959(.A(n1000), .O(n999));
  andx g0960(.A(pi05), .B(pi18), .O(n1000));
  andx g0961(.A(pi00), .B(pi07), .O(n1001));
  orx  g0962(.A(n1006), .B(n1003), .O(n1002));
  invx g0963(.A(n1004), .O(n1003));
  orx  g0964(.A(n1005), .B(n1007), .O(n1004));
  andx g0965(.A(pi15), .B(pi10), .O(n1005));
  andx g0966(.A(n1007), .B(pi10), .O(n1006));
  orx  g0967(.A(n1009), .B(n1008), .O(n1007));
  andx g0968(.A(n1096), .B(n1097), .O(n1008));
  andx g0969(.A(n1092), .B(n1010), .O(n1009));
  orx  g0970(.A(n1096), .B(n1097), .O(n1010));
  orx  g0971(.A(n1013), .B(n1012), .O(n1011));
  andx g0972(.A(n1016), .B(pi13), .O(n1012));
  andx g0973(.A(n1015), .B(n1014), .O(n1013));
  orx  g0974(.A(n1117), .B(n1149), .O(n1014));
  invx g0975(.A(n1016), .O(n1015));
  orx  g0976(.A(n1017), .B(n1108), .O(n1016));
  andx g0977(.A(n1085), .B(n1106), .O(n1017));
  orx  g0978(.A(n1022), .B(n1019), .O(n1018));
  invx g0979(.A(n1020), .O(n1019));
  orx  g0980(.A(n1021), .B(n1023), .O(n1020));
  andx g0981(.A(pi14), .B(pi11), .O(n1021));
  andx g0982(.A(n1023), .B(pi14), .O(n1022));
  orx  g0983(.A(n1024), .B(n1114), .O(n1023));
  andx g0984(.A(n1081), .B(n1025), .O(n1024));
  orx  g0985(.A(n1026), .B(n1119), .O(n1025));
  andx g0986(.A(pi13), .B(pi11), .O(n1026));
  orx  g0987(.A(n1029), .B(n1028), .O(n1027));
  andx g0988(.A(n1033), .B(pi16), .O(n1028));
  andx g0989(.A(n1032), .B(n1030), .O(n1029));
  orx  g0990(.A(n1059), .B(n1031), .O(n1030));
  invx g0991(.A(pi16), .O(n1031));
  invx g0992(.A(n1033), .O(n1032));
  orx  g0993(.A(n1035), .B(n1034), .O(n1033));
  andx g0994(.A(n1037), .B(pi14), .O(n1034));
  andx g0995(.A(n1077), .B(n1036), .O(n1035));
  orx  g0996(.A(n1076), .B(n1037), .O(n1036));
  orx  g0997(.A(n1039), .B(n1038), .O(n1037));
  andx g0998(.A(n1041), .B(pi13), .O(n1038));
  andx g0999(.A(n1070), .B(n1040), .O(n1039));
  orx  g1000(.A(n1069), .B(n1041), .O(n1040));
  orx  g1001(.A(n1043), .B(n1042), .O(n1041));
  andx g1002(.A(n1045), .B(pi10), .O(n1042));
  andx g1003(.A(n1061), .B(n1044), .O(n1043));
  orx  g1004(.A(n1060), .B(n1045), .O(n1044));
  orx  g1005(.A(n1047), .B(n1046), .O(n1045));
  andx g1006(.A(n1055), .B(n1049), .O(n1046));
  andx g1007(.A(n1056), .B(n1048), .O(n1047));
  orx  g1008(.A(n1055), .B(n1049), .O(n1048));
  orx  g1009(.A(n1051), .B(n1050), .O(n1049));
  andx g1010(.A(n1053), .B(n1054), .O(n1050));
  invx g1011(.A(n1052), .O(n1051));
  orx  g1012(.A(n1054), .B(n1053), .O(n1052));
  andx g1013(.A(pi00), .B(pi12), .O(n1053));
  orx  g1014(.A(n1161), .B(n1137), .O(n1054));
  andx g1015(.A(pi08), .B(pi09), .O(n1055));
  invx g1016(.A(n1057), .O(n1056));
  orx  g1017(.A(n41), .B(n1058), .O(n1057));
  orx  g1018(.A(n1059), .B(n1137), .O(n1058));
  invx g1019(.A(pi09), .O(n1059));
  andx g1020(.A(pi10), .B(pi09), .O(n1060));
  orx  g1021(.A(n1064), .B(n1062), .O(n1061));
  invx g1022(.A(n1063), .O(n1062));
  orx  g1023(.A(n1065), .B(n1127), .O(n1063));
  andx g1024(.A(n1127), .B(n1065), .O(n1064));
  andx g1025(.A(n1067), .B(n1066), .O(n1065));
  orx  g1026(.A(n1135), .B(n1133), .O(n1066));
  orx  g1027(.A(n1068), .B(n1134), .O(n1067));
  invx g1028(.A(n1133), .O(n1068));
  andx g1029(.A(pi13), .B(pi09), .O(n1069));
  orx  g1030(.A(n1072), .B(n1071), .O(n1070));
  andx g1031(.A(n1139), .B(n1074), .O(n1071));
  invx g1032(.A(n1073), .O(n1072));
  orx  g1033(.A(n1074), .B(n1139), .O(n1073));
  orx  g1034(.A(n1120), .B(n1075), .O(n1074));
  invx g1035(.A(n1122), .O(n1075));
  andx g1036(.A(pi14), .B(pi09), .O(n1076));
  orx  g1037(.A(n1079), .B(n1078), .O(n1077));
  andx g1038(.A(n1081), .B(n1113), .O(n1078));
  invx g1039(.A(n1080), .O(n1079));
  orx  g1040(.A(n1113), .B(n1081), .O(n1080));
  orx  g1041(.A(n1083), .B(n1082), .O(n1081));
  andx g1042(.A(n1085), .B(n1104), .O(n1082));
  invx g1043(.A(n1084), .O(n1083));
  orx  g1044(.A(n1104), .B(n1085), .O(n1084));
  orx  g1045(.A(n1088), .B(n1086), .O(n1085));
  invx g1046(.A(n1087), .O(n1086));
  orx  g1047(.A(n1089), .B(n1097), .O(n1087));
  andx g1048(.A(n1097), .B(n1089), .O(n1088));
  andx g1049(.A(n1091), .B(n1090), .O(n1089));
  orx  g1050(.A(n1093), .B(n1096), .O(n1090));
  orx  g1051(.A(n1095), .B(n1092), .O(n1091));
  invx g1052(.A(n1093), .O(n1092));
  orx  g1053(.A(n1103), .B(n1094), .O(n1093));
  orx  g1054(.A(n41), .B(n1160), .O(n1094));
  invx g1055(.A(n1096), .O(n1095));
  andx g1056(.A(pi08), .B(pi15), .O(n1096));
  orx  g1057(.A(n1099), .B(n1098), .O(n1097));
  andx g1058(.A(n1101), .B(n1102), .O(n1098));
  invx g1059(.A(n1100), .O(n1099));
  orx  g1060(.A(n1102), .B(n1101), .O(n1100));
  andx g1061(.A(pi00), .B(pi18), .O(n1101));
  orx  g1062(.A(n1161), .B(n1103), .O(n1102));
  invx g1063(.A(pi17), .O(n1103));
  orx  g1064(.A(n1108), .B(n1105), .O(n1104));
  invx g1065(.A(n1106), .O(n1105));
  orx  g1066(.A(n1107), .B(n1109), .O(n1106));
  andx g1067(.A(pi12), .B(pi10), .O(n1107));
  andx g1068(.A(n1109), .B(pi10), .O(n1108));
  orx  g1069(.A(n1111), .B(n1110), .O(n1109));
  andx g1070(.A(n1153), .B(n1154), .O(n1110));
  andx g1071(.A(n1146), .B(n1112), .O(n1111));
  orx  g1072(.A(n1153), .B(n1154), .O(n1112));
  orx  g1073(.A(n1115), .B(n1114), .O(n1113));
  andx g1074(.A(n1119), .B(pi13), .O(n1114));
  andx g1075(.A(n1118), .B(n1116), .O(n1115));
  orx  g1076(.A(n1137), .B(n1117), .O(n1116));
  invx g1077(.A(pi13), .O(n1117));
  invx g1078(.A(n1119), .O(n1118));
  orx  g1079(.A(n1121), .B(n1120), .O(n1119));
  andx g1080(.A(n1123), .B(pi10), .O(n1120));
  andx g1081(.A(n1139), .B(n1122), .O(n1121));
  orx  g1082(.A(n1138), .B(n1123), .O(n1122));
  orx  g1083(.A(n1125), .B(n1124), .O(n1123));
  andx g1084(.A(n1133), .B(n1127), .O(n1124));
  andx g1085(.A(n1134), .B(n1126), .O(n1125));
  orx  g1086(.A(n1133), .B(n1127), .O(n1126));
  orx  g1087(.A(n1129), .B(n1128), .O(n1127));
  andx g1088(.A(n1131), .B(n1132), .O(n1128));
  invx g1089(.A(n1130), .O(n1129));
  orx  g1090(.A(n1132), .B(n1131), .O(n1130));
  andx g1091(.A(pi00), .B(pi15), .O(n1131));
  orx  g1092(.A(n1161), .B(n1149), .O(n1132));
  andx g1093(.A(pi08), .B(pi11), .O(n1133));
  invx g1094(.A(n1135), .O(n1134));
  orx  g1095(.A(n1149), .B(n1136), .O(n1135));
  orx  g1096(.A(n1137), .B(n41), .O(n1136));
  invx g1097(.A(pi11), .O(n1137));
  andx g1098(.A(pi11), .B(pi10), .O(n1138));
  orx  g1099(.A(n1142), .B(n1140), .O(n1139));
  invx g1100(.A(n1141), .O(n1140));
  orx  g1101(.A(n1143), .B(n1154), .O(n1141));
  andx g1102(.A(n1154), .B(n1143), .O(n1142));
  andx g1103(.A(n1145), .B(n1144), .O(n1143));
  orx  g1104(.A(n1147), .B(n1153), .O(n1144));
  orx  g1105(.A(n1152), .B(n1146), .O(n1145));
  invx g1106(.A(n1147), .O(n1146));
  orx  g1107(.A(n1160), .B(n1148), .O(n1147));
  orx  g1108(.A(n41), .B(n1149), .O(n1148));
  invx g1109(.A(pi12), .O(n1149));
  orx  g1110(.A(n1151), .B(n40), .O(n1150));
  invx g1111(.A(pi00), .O(n1151));
  invx g1112(.A(n1153), .O(n1152));
  andx g1113(.A(pi08), .B(pi12), .O(n1153));
  orx  g1114(.A(n1156), .B(n1155), .O(n1154));
  andx g1115(.A(n1158), .B(n1159), .O(n1155));
  invx g1116(.A(n1157), .O(n1156));
  orx  g1117(.A(n1159), .B(n1158), .O(n1157));
  andx g1118(.A(pi00), .B(pi17), .O(n1158));
  orx  g1119(.A(n1161), .B(n1160), .O(n1159));
  invx g1120(.A(pi15), .O(n1160));
  invx g1121(.A(pi05), .O(n1161));
  andx g1122(.A(pi00), .B(pi01), .O(po00));
endmodule


