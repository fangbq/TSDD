// Benchmark "top" written by ABC on Fri Feb  7 13:36:32 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13;
  wire n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
    n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
    n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
    n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
    n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
    n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294;
  invx g0000(.a(pi09), .O(n28));
  invx g0001(.a(pi13), .O(n29));
  andx g0002(.a(n29), .b(pi12), .O(n30));
  andx g0003(.a(n30), .b(n28), .O(n31));
  andx g0004(.a(pi10), .b(pi08), .O(n32));
  andx g0005(.a(n32), .b(n31), .O(n33));
  andx g0006(.a(pi03), .b(pi01), .O(n34));
  andx g0007(.a(n34), .b(pi00), .O(n35));
  invx g0008(.a(pi02), .O(n36));
  invx g0009(.a(pi04), .O(n37));
  andx g0010(.a(pi06), .b(n37), .O(n38));
  andx g0011(.a(n38), .b(n36), .O(n39));
  andx g0012(.a(n39), .b(n35), .O(n40));
  invx g0013(.a(pi05), .O(n41));
  andx g0014(.a(pi06), .b(n41), .O(n42));
  andx g0015(.a(n42), .b(n37), .O(n43));
  andx g0016(.a(n43), .b(n35), .O(n44));
  orx  g0017(.a(n44), .b(n40), .O(n45));
  andx g0018(.a(n45), .b(n33), .O(n46));
  andx g0019(.a(n35), .b(n29), .O(n47));
  invx g0020(.a(pi06), .O(n48));
  andx g0021(.a(n37), .b(pi03), .O(n49));
  andx g0022(.a(n49), .b(n48), .O(n50));
  andx g0023(.a(pi12), .b(pi10), .O(n51));
  andx g0024(.a(n51), .b(pi07), .O(n52));
  andx g0025(.a(n52), .b(n50), .O(n53));
  andx g0026(.a(n53), .b(n47), .O(n54));
  orx  g0027(.a(n54), .b(n46), .O(n55));
  andx g0028(.a(n36), .b(pi01), .O(n56));
  andx g0029(.a(n56), .b(pi00), .O(n57));
  andx g0030(.a(n57), .b(n50), .O(n58));
  invx g0031(.a(pi03), .O(n59));
  andx g0032(.a(pi02), .b(pi01), .O(n60));
  andx g0033(.a(n60), .b(pi00), .O(n61));
  andx g0034(.a(n61), .b(n59), .O(n62));
  andx g0035(.a(pi04), .b(pi02), .O(n63));
  andx g0036(.a(n63), .b(n48), .O(n64));
  andx g0037(.a(n64), .b(n62), .O(n65));
  orx  g0038(.a(n65), .b(n58), .O(n66));
  andx g0039(.a(pi10), .b(pi07), .O(n67));
  andx g0040(.a(n67), .b(n48), .O(n68));
  andx g0041(.a(n68), .b(n30), .O(n69));
  andx g0042(.a(n69), .b(n66), .O(n70));
  invx g0043(.a(pi08), .O(n71));
  andx g0044(.a(n71), .b(pi07), .O(n72));
  invx g0045(.a(pi12), .O(n73));
  andx g0046(.a(n29), .b(n73), .O(n74));
  andx g0047(.a(n74), .b(n72), .O(n75));
  andx g0048(.a(n75), .b(pi10), .O(n76));
  invx g0049(.a(pi07), .O(n77));
  andx g0050(.a(n32), .b(n77), .O(n78));
  andx g0051(.a(n78), .b(n74), .O(n79));
  orx  g0052(.a(n79), .b(n76), .O(n80));
  invx g0053(.a(pi10), .O(n81));
  andx g0054(.a(n81), .b(pi09), .O(n82));
  andx g0055(.a(n82), .b(pi07), .O(n83));
  andx g0056(.a(n83), .b(n74), .O(n84));
  andx g0057(.a(n74), .b(n28), .O(n85));
  andx g0058(.a(n85), .b(n67), .O(n86));
  orx  g0059(.a(n86), .b(n84), .O(n87));
  orx  g0060(.a(n87), .b(n80), .O(n88));
  andx g0061(.a(pi04), .b(pi03), .O(n89));
  andx g0062(.a(n89), .b(pi02), .O(n90));
  andx g0063(.a(n90), .b(n41), .O(n91));
  andx g0064(.a(n91), .b(n88), .O(n92));
  orx  g0065(.a(n92), .b(n70), .O(n93));
  orx  g0066(.a(n93), .b(n55), .O(n94));
  andx g0067(.a(n63), .b(pi01), .O(n95));
  andx g0068(.a(pi07), .b(n41), .O(n96));
  andx g0069(.a(n96), .b(n59), .O(n97));
  andx g0070(.a(n97), .b(n95), .O(n98));
  invx g0071(.a(pi11), .O(n99));
  andx g0072(.a(pi13), .b(n73), .O(n100));
  andx g0073(.a(n100), .b(n99), .O(n101));
  andx g0074(.a(n101), .b(n67), .O(n102));
  andx g0075(.a(n100), .b(pi10), .O(n103));
  andx g0076(.a(n103), .b(n71), .O(n104));
  orx  g0077(.a(n104), .b(n102), .O(n105));
  andx g0078(.a(n105), .b(n98), .O(n106));
  andx g0079(.a(n95), .b(pi13), .O(n107));
  andx g0080(.a(pi07), .b(pi06), .O(n108));
  andx g0081(.a(n108), .b(n41), .O(n109));
  andx g0082(.a(n73), .b(pi10), .O(n110));
  andx g0083(.a(n110), .b(n71), .O(n111));
  andx g0084(.a(n111), .b(n109), .O(n112));
  andx g0085(.a(n73), .b(n99), .O(n113));
  andx g0086(.a(n113), .b(pi10), .O(n114));
  andx g0087(.a(n114), .b(n109), .O(n115));
  orx  g0088(.a(n115), .b(n112), .O(n116));
  andx g0089(.a(n116), .b(n107), .O(n117));
  orx  g0090(.a(n117), .b(n106), .O(n118));
  andx g0091(.a(n30), .b(n99), .O(n119));
  andx g0092(.a(pi09), .b(pi07), .O(n120));
  andx g0093(.a(n120), .b(n119), .O(n121));
  andx g0094(.a(n82), .b(n71), .O(n122));
  andx g0095(.a(n122), .b(n30), .O(n123));
  orx  g0096(.a(n123), .b(n121), .O(n124));
  andx g0097(.a(n124), .b(n40), .O(n125));
  andx g0098(.a(n38), .b(n35), .O(n126));
  andx g0099(.a(n126), .b(n121), .O(n127));
  orx  g0100(.a(n127), .b(n125), .O(n128));
  orx  g0101(.a(n128), .b(n118), .O(n129));
  andx g0102(.a(pi11), .b(n28), .O(n130));
  andx g0103(.a(n30), .b(pi07), .O(n131));
  andx g0104(.a(n131), .b(n130), .O(n132));
  andx g0105(.a(n48), .b(n41), .O(n133));
  andx g0106(.a(n133), .b(n37), .O(n134));
  andx g0107(.a(n134), .b(n35), .O(n135));
  orx  g0108(.a(n135), .b(n65), .O(n136));
  andx g0109(.a(n136), .b(n132), .O(n137));
  andx g0110(.a(pi04), .b(n59), .O(n138));
  andx g0111(.a(n138), .b(pi01), .O(n139));
  andx g0112(.a(n139), .b(n29), .O(n140));
  andx g0113(.a(pi08), .b(pi06), .O(n141));
  andx g0114(.a(n141), .b(n41), .O(n142));
  andx g0115(.a(n51), .b(n28), .O(n143));
  andx g0116(.a(n143), .b(n142), .O(n144));
  andx g0117(.a(pi12), .b(n99), .O(n145));
  andx g0118(.a(n145), .b(pi10), .O(n146));
  andx g0119(.a(n28), .b(pi06), .O(n147));
  andx g0120(.a(n147), .b(n41), .O(n148));
  andx g0121(.a(n148), .b(n146), .O(n149));
  orx  g0122(.a(n149), .b(n144), .O(n150));
  andx g0123(.a(n71), .b(pi06), .O(n151));
  andx g0124(.a(n151), .b(n41), .O(n152));
  andx g0125(.a(pi12), .b(pi11), .O(n153));
  andx g0126(.a(n153), .b(pi09), .O(n154));
  andx g0127(.a(n154), .b(n152), .O(n155));
  andx g0128(.a(n146), .b(n142), .O(n156));
  orx  g0129(.a(n156), .b(n155), .O(n157));
  orx  g0130(.a(n157), .b(n150), .O(n158));
  andx g0131(.a(n158), .b(n140), .O(n159));
  orx  g0132(.a(n159), .b(n137), .O(n160));
  orx  g0133(.a(n160), .b(n129), .O(n161));
  andx g0134(.a(n30), .b(n81), .O(n162));
  andx g0135(.a(pi11), .b(pi09), .O(n163));
  andx g0136(.a(n163), .b(n162), .O(n164));
  andx g0137(.a(n164), .b(n40), .O(n165));
  invx g0138(.a(n89), .O(n166));
  andx g0139(.a(pi05), .b(pi02), .O(n167));
  andx g0140(.a(n167), .b(n166), .O(n168));
  andx g0141(.a(n168), .b(n76), .O(n169));
  orx  g0142(.a(n169), .b(n165), .O(n170));
  andx g0143(.a(n99), .b(pi10), .O(n171));
  andx g0144(.a(n171), .b(n31), .O(n172));
  andx g0145(.a(pi06), .b(pi04), .O(n173));
  andx g0146(.a(n173), .b(n59), .O(n174));
  andx g0147(.a(n174), .b(n61), .O(n175));
  andx g0148(.a(n175), .b(n172), .O(n176));
  andx g0149(.a(n59), .b(pi02), .O(n177));
  andx g0150(.a(n177), .b(pi01), .O(n178));
  andx g0151(.a(n178), .b(pi13), .O(n179));
  andx g0152(.a(n77), .b(pi06), .O(n180));
  andx g0153(.a(n180), .b(n37), .O(n181));
  andx g0154(.a(n110), .b(pi08), .O(n182));
  andx g0155(.a(n182), .b(n181), .O(n183));
  andx g0156(.a(n183), .b(n179), .O(n184));
  orx  g0157(.a(n184), .b(n176), .O(n185));
  orx  g0158(.a(n185), .b(n170), .O(n186));
  andx g0159(.a(pi05), .b(n37), .O(n187));
  andx g0160(.a(n187), .b(pi02), .O(n188));
  andx g0161(.a(n188), .b(n86), .O(n189));
  andx g0162(.a(pi05), .b(pi04), .O(n190));
  andx g0163(.a(n190), .b(n59), .O(n191));
  andx g0164(.a(n191), .b(n57), .O(n192));
  andx g0165(.a(n30), .b(pi11), .O(n193));
  andx g0166(.a(n82), .b(pi06), .O(n194));
  andx g0167(.a(n194), .b(n193), .O(n195));
  andx g0168(.a(n195), .b(n192), .O(n196));
  orx  g0169(.a(n196), .b(n189), .O(n197));
  andx g0170(.a(pi05), .b(n59), .O(n198));
  andx g0171(.a(n198), .b(pi02), .O(n199));
  andx g0172(.a(n199), .b(n84), .O(n200));
  andx g0173(.a(pi08), .b(n77), .O(n201));
  andx g0174(.a(n201), .b(pi11), .O(n202));
  andx g0175(.a(n202), .b(n30), .O(n203));
  andx g0176(.a(n203), .b(n40), .O(n204));
  orx  g0177(.a(n204), .b(n200), .O(n205));
  orx  g0178(.a(n205), .b(n197), .O(n206));
  orx  g0179(.a(n206), .b(n186), .O(n207));
  andx g0180(.a(n130), .b(pi08), .O(n208));
  andx g0181(.a(n180), .b(pi05), .O(n209));
  andx g0182(.a(n209), .b(n208), .O(n210));
  andx g0183(.a(n139), .b(n100), .O(n211));
  andx g0184(.a(n211), .b(n210), .O(n212));
  andx g0185(.a(n77), .b(n41), .O(n213));
  andx g0186(.a(n213), .b(pi04), .O(n214));
  andx g0187(.a(n214), .b(n178), .O(n215));
  andx g0188(.a(n100), .b(pi08), .O(n216));
  andx g0189(.a(n216), .b(n130), .O(n217));
  andx g0190(.a(n217), .b(n215), .O(n218));
  orx  g0191(.a(n218), .b(n212), .O(n219));
  andx g0192(.a(n67), .b(n49), .O(n220));
  andx g0193(.a(n220), .b(n119), .O(n221));
  andx g0194(.a(n221), .b(n57), .O(n222));
  andx g0195(.a(n67), .b(pi04), .O(n223));
  andx g0196(.a(n223), .b(n119), .O(n224));
  andx g0197(.a(n224), .b(n62), .O(n225));
  orx  g0198(.a(n225), .b(n222), .O(n226));
  orx  g0199(.a(n226), .b(n219), .O(n227));
  andx g0200(.a(n35), .b(n30), .O(n228));
  andx g0201(.a(pi06), .b(pi05), .O(n229));
  andx g0202(.a(n229), .b(n37), .O(n230));
  andx g0203(.a(n171), .b(pi08), .O(n231));
  andx g0204(.a(n231), .b(n230), .O(n232));
  andx g0205(.a(n232), .b(n228), .O(n233));
  andx g0206(.a(n145), .b(pi09), .O(n234));
  andx g0207(.a(n234), .b(n109), .O(n235));
  andx g0208(.a(n235), .b(n140), .O(n236));
  orx  g0209(.a(n236), .b(n233), .O(n237));
  andx g0210(.a(n172), .b(n40), .O(n238));
  andx g0211(.a(n139), .b(pi13), .O(n239));
  andx g0212(.a(n108), .b(pi05), .O(n240));
  andx g0213(.a(n73), .b(n81), .O(n241));
  andx g0214(.a(n241), .b(pi09), .O(n242));
  andx g0215(.a(n242), .b(n240), .O(n243));
  andx g0216(.a(n243), .b(n239), .O(n244));
  orx  g0217(.a(n244), .b(n238), .O(n245));
  orx  g0218(.a(n245), .b(n237), .O(n246));
  orx  g0219(.a(n246), .b(n227), .O(n247));
  orx  g0220(.a(n247), .b(n207), .O(n248));
  orx  g0221(.a(n248), .b(n161), .O(n249));
  orx  g0222(.a(n249), .b(n94), .O(n250));
  orx  g0223(.a(n175), .b(n44), .O(n251));
  andx g0224(.a(n251), .b(n203), .O(n252));
  andx g0225(.a(pi03), .b(n36), .O(n253));
  andx g0226(.a(n253), .b(pi01), .O(n254));
  andx g0227(.a(pi07), .b(n48), .O(n255));
  andx g0228(.a(n255), .b(pi05), .O(n256));
  andx g0229(.a(n256), .b(n254), .O(n257));
  andx g0230(.a(n255), .b(n41), .O(n258));
  andx g0231(.a(n258), .b(n95), .O(n259));
  orx  g0232(.a(n259), .b(n257), .O(n260));
  andx g0233(.a(n260), .b(n105), .O(n261));
  orx  g0234(.a(n261), .b(n252), .O(n262));
  andx g0235(.a(n251), .b(n164), .O(n263));
  andx g0236(.a(n67), .b(pi05), .O(n264));
  andx g0237(.a(n264), .b(n119), .O(n265));
  andx g0238(.a(n30), .b(pi10), .O(n266));
  andx g0239(.a(n266), .b(n256), .O(n267));
  orx  g0240(.a(n267), .b(n265), .O(n268));
  andx g0241(.a(n268), .b(n192), .O(n269));
  orx  g0242(.a(n269), .b(n263), .O(n270));
  orx  g0243(.a(n270), .b(n262), .O(n271));
  andx g0244(.a(n153), .b(n28), .O(n272));
  andx g0245(.a(n272), .b(n258), .O(n273));
  andx g0246(.a(n273), .b(n140), .O(n274));
  andx g0247(.a(pi04), .b(pi01), .O(n275));
  invx g0248(.a(pi00), .O(n276));
  andx g0249(.a(n29), .b(n276), .O(n277));
  andx g0250(.a(n277), .b(n275), .O(n278));
  andx g0251(.a(n171), .b(n30), .O(n279));
  andx g0252(.a(n279), .b(pi07), .O(n280));
  andx g0253(.a(n280), .b(n278), .O(n281));
  orx  g0254(.a(n281), .b(n274), .O(n282));
  andx g0255(.a(n110), .b(n28), .O(n283));
  andx g0256(.a(n283), .b(n240), .O(n284));
  andx g0257(.a(n284), .b(n239), .O(n285));
  andx g0258(.a(n56), .b(pi13), .O(n286));
  andx g0259(.a(n286), .b(pi03), .O(n287));
  andx g0260(.a(n287), .b(n243), .O(n288));
  orx  g0261(.a(n288), .b(n285), .O(n289));
  orx  g0262(.a(n289), .b(n282), .O(n290));
  andx g0263(.a(n67), .b(n41), .O(n291));
  andx g0264(.a(n291), .b(n119), .O(n292));
  andx g0265(.a(n153), .b(n42), .O(n293));
  andx g0266(.a(n293), .b(n82), .O(n294));
  orx  g0267(.a(n294), .b(n292), .O(n295));
  andx g0268(.a(n295), .b(n140), .O(n296));
  andx g0269(.a(n74), .b(n99), .O(n297));
  andx g0270(.a(n297), .b(n67), .O(n298));
  andx g0271(.a(n298), .b(n91), .O(n299));
  andx g0272(.a(n90), .b(n29), .O(n300));
  andx g0273(.a(n73), .b(pi11), .O(n301));
  andx g0274(.a(n301), .b(n28), .O(n302));
  andx g0275(.a(n201), .b(n41), .O(n303));
  andx g0276(.a(n303), .b(n302), .O(n304));
  andx g0277(.a(n304), .b(n300), .O(n305));
  orx  g0278(.a(n305), .b(n299), .O(n306));
  orx  g0279(.a(n306), .b(n296), .O(n307));
  orx  g0280(.a(n307), .b(n290), .O(n308));
  orx  g0281(.a(n308), .b(n271), .O(n309));
  andx g0282(.a(n187), .b(pi01), .O(n310));
  andx g0283(.a(n201), .b(n48), .O(n311));
  andx g0284(.a(n311), .b(n103), .O(n312));
  andx g0285(.a(n312), .b(n310), .O(n313));
  andx g0286(.a(n49), .b(pi01), .O(n314));
  andx g0287(.a(n201), .b(pi05), .O(n315));
  andx g0288(.a(n315), .b(n103), .O(n316));
  andx g0289(.a(n316), .b(n314), .O(n317));
  orx  g0290(.a(n317), .b(n313), .O(n318));
  andx g0291(.a(n209), .b(n182), .O(n319));
  orx  g0292(.a(n287), .b(n239), .O(n320));
  andx g0293(.a(n320), .b(n319), .O(n321));
  orx  g0294(.a(n321), .b(n318), .O(n322));
  andx g0295(.a(n275), .b(n276), .O(n323));
  andx g0296(.a(n323), .b(n69), .O(n324));
  andx g0297(.a(n199), .b(n79), .O(n325));
  orx  g0298(.a(n325), .b(n324), .O(n326));
  andx g0299(.a(pi09), .b(n71), .O(n327));
  andx g0300(.a(n327), .b(pi06), .O(n328));
  andx g0301(.a(n328), .b(n192), .O(n329));
  andx g0302(.a(n329), .b(n193), .O(n330));
  orx  g0303(.a(n330), .b(n326), .O(n331));
  orx  g0304(.a(n331), .b(n322), .O(n332));
  andx g0305(.a(n279), .b(n141), .O(n333));
  andx g0306(.a(n279), .b(n147), .O(n334));
  orx  g0307(.a(n334), .b(n333), .O(n335));
  andx g0308(.a(n335), .b(n192), .O(n336));
  andx g0309(.a(n230), .b(n202), .O(n337));
  andx g0310(.a(n337), .b(n228), .O(n338));
  andx g0311(.a(n72), .b(pi11), .O(n339));
  andx g0312(.a(n339), .b(n30), .O(n340));
  andx g0313(.a(n340), .b(n40), .O(n341));
  orx  g0314(.a(n341), .b(n338), .O(n342));
  orx  g0315(.a(n342), .b(n336), .O(n343));
  andx g0316(.a(n231), .b(n30), .O(n344));
  orx  g0317(.a(n344), .b(n123), .O(n345));
  andx g0318(.a(n345), .b(n251), .O(n346));
  andx g0319(.a(n72), .b(n48), .O(n347));
  andx g0320(.a(n347), .b(n103), .O(n348));
  andx g0321(.a(n348), .b(n310), .O(n349));
  andx g0322(.a(n72), .b(pi05), .O(n350));
  andx g0323(.a(n314), .b(n103), .O(n351));
  andx g0324(.a(n351), .b(n350), .O(n352));
  orx  g0325(.a(n352), .b(n349), .O(n353));
  orx  g0326(.a(n353), .b(n346), .O(n354));
  orx  g0327(.a(n354), .b(n343), .O(n355));
  orx  g0328(.a(n355), .b(n332), .O(n356));
  orx  g0329(.a(n356), .b(n309), .O(n357));
  andx g0330(.a(n108), .b(n37), .O(n358));
  andx g0331(.a(n358), .b(n111), .O(n359));
  andx g0332(.a(n359), .b(n179), .O(n360));
  andx g0333(.a(n180), .b(n41), .O(n361));
  andx g0334(.a(n153), .b(pi08), .O(n362));
  andx g0335(.a(n362), .b(n361), .O(n363));
  andx g0336(.a(n363), .b(n140), .O(n364));
  orx  g0337(.a(n364), .b(n360), .O(n365));
  andx g0338(.a(n334), .b(n323), .O(n366));
  andx g0339(.a(n323), .b(n195), .O(n367));
  orx  g0340(.a(n367), .b(n366), .O(n368));
  orx  g0341(.a(n368), .b(n365), .O(n369));
  andx g0342(.a(n358), .b(n114), .O(n370));
  andx g0343(.a(n370), .b(n179), .O(n371));
  andx g0344(.a(n361), .b(n182), .O(n372));
  andx g0345(.a(n372), .b(n107), .O(n373));
  orx  g0346(.a(n373), .b(n371), .O(n374));
  andx g0347(.a(n240), .b(n114), .O(n375));
  andx g0348(.a(n375), .b(n287), .O(n376));
  andx g0349(.a(n221), .b(n35), .O(n377));
  orx  g0350(.a(n377), .b(n376), .O(n378));
  orx  g0351(.a(n378), .b(n374), .O(n379));
  orx  g0352(.a(n379), .b(n369), .O(n380));
  andx g0353(.a(pi11), .b(n81), .O(n381));
  andx g0354(.a(n381), .b(pi09), .O(n382));
  andx g0355(.a(n382), .b(n230), .O(n383));
  andx g0356(.a(n383), .b(n228), .O(n384));
  andx g0357(.a(n77), .b(n48), .O(n385));
  andx g0358(.a(n385), .b(pi05), .O(n386));
  andx g0359(.a(n386), .b(n254), .O(n387));
  andx g0360(.a(n387), .b(n217), .O(n388));
  orx  g0361(.a(n388), .b(n384), .O(n389));
  andx g0362(.a(n208), .b(n181), .O(n390));
  andx g0363(.a(n178), .b(n100), .O(n391));
  andx g0364(.a(n391), .b(n390), .O(n392));
  andx g0365(.a(n254), .b(n100), .O(n393));
  andx g0366(.a(n393), .b(n210), .O(n394));
  orx  g0367(.a(n394), .b(n392), .O(n395));
  orx  g0368(.a(n395), .b(n389), .O(n396));
  andx g0369(.a(n28), .b(pi07), .O(n397));
  andx g0370(.a(n397), .b(pi05), .O(n398));
  andx g0371(.a(n398), .b(n314), .O(n399));
  andx g0372(.a(n399), .b(n103), .O(n400));
  andx g0373(.a(n397), .b(n48), .O(n401));
  andx g0374(.a(n401), .b(n103), .O(n402));
  andx g0375(.a(n402), .b(n310), .O(n403));
  orx  g0376(.a(n403), .b(n400), .O(n404));
  andx g0377(.a(n199), .b(n86), .O(n405));
  andx g0378(.a(n201), .b(pi06), .O(n406));
  andx g0379(.a(n406), .b(n193), .O(n407));
  andx g0380(.a(n407), .b(n192), .O(n408));
  orx  g0381(.a(n408), .b(n405), .O(n409));
  orx  g0382(.a(n409), .b(n404), .O(n410));
  orx  g0383(.a(n410), .b(n396), .O(n411));
  orx  g0384(.a(n411), .b(n380), .O(n412));
  andx g0385(.a(n101), .b(n68), .O(n413));
  andx g0386(.a(n413), .b(n310), .O(n414));
  andx g0387(.a(n240), .b(n111), .O(n415));
  andx g0388(.a(n415), .b(n239), .O(n416));
  orx  g0389(.a(n416), .b(n414), .O(n417));
  andx g0390(.a(n340), .b(n126), .O(n418));
  andx g0391(.a(n28), .b(pi08), .O(n419));
  andx g0392(.a(n419), .b(n77), .O(n420));
  andx g0393(.a(n74), .b(pi11), .O(n421));
  andx g0394(.a(n421), .b(n420), .O(n422));
  andx g0395(.a(n422), .b(n168), .O(n423));
  orx  g0396(.a(n423), .b(n418), .O(n424));
  orx  g0397(.a(n424), .b(n417), .O(n425));
  andx g0398(.a(n358), .b(n242), .O(n426));
  andx g0399(.a(n426), .b(n179), .O(n427));
  andx g0400(.a(n264), .b(n101), .O(n428));
  andx g0401(.a(n428), .b(n314), .O(n429));
  orx  g0402(.a(n429), .b(n427), .O(n430));
  andx g0403(.a(n358), .b(n283), .O(n431));
  andx g0404(.a(n431), .b(n179), .O(n432));
  andx g0405(.a(n287), .b(n284), .O(n433));
  orx  g0406(.a(n433), .b(n432), .O(n434));
  orx  g0407(.a(n434), .b(n430), .O(n435));
  orx  g0408(.a(n435), .b(n425), .O(n436));
  andx g0409(.a(n175), .b(n121), .O(n437));
  andx g0410(.a(n48), .b(pi05), .O(n438));
  andx g0411(.a(n438), .b(n37), .O(n439));
  andx g0412(.a(n130), .b(pi07), .O(n440));
  andx g0413(.a(n440), .b(n439), .O(n441));
  andx g0414(.a(n441), .b(n228), .O(n442));
  orx  g0415(.a(n442), .b(n437), .O(n443));
  andx g0416(.a(n188), .b(n84), .O(n444));
  andx g0417(.a(n298), .b(n199), .O(n445));
  orx  g0418(.a(n445), .b(n444), .O(n446));
  orx  g0419(.a(n446), .b(n443), .O(n447));
  andx g0420(.a(n340), .b(n175), .O(n448));
  andx g0421(.a(n132), .b(n58), .O(n449));
  orx  g0422(.a(n449), .b(n448), .O(n450));
  andx g0423(.a(n415), .b(n287), .O(n451));
  andx g0424(.a(n182), .b(pi13), .O(n452));
  andx g0425(.a(n452), .b(n215), .O(n453));
  orx  g0426(.a(n453), .b(n451), .O(n454));
  orx  g0427(.a(n454), .b(n450), .O(n455));
  orx  g0428(.a(n455), .b(n447), .O(n456));
  orx  g0429(.a(n456), .b(n436), .O(n457));
  orx  g0430(.a(n457), .b(n412), .O(n458));
  orx  g0431(.a(n458), .b(n357), .O(n459));
  andx g0432(.a(n401), .b(n193), .O(n460));
  andx g0433(.a(n340), .b(pi06), .O(n461));
  orx  g0434(.a(n461), .b(n460), .O(n462));
  andx g0435(.a(n328), .b(n162), .O(n463));
  andx g0436(.a(n328), .b(n193), .O(n464));
  orx  g0437(.a(n464), .b(n463), .O(n465));
  andx g0438(.a(n120), .b(pi06), .O(n466));
  andx g0439(.a(n466), .b(n119), .O(n467));
  orx  g0440(.a(n467), .b(n407), .O(n468));
  orx  g0441(.a(n468), .b(n465), .O(n469));
  orx  g0442(.a(n469), .b(n462), .O(n470));
  andx g0443(.a(n470), .b(n323), .O(n471));
  andx g0444(.a(n419), .b(pi06), .O(n472));
  andx g0445(.a(n472), .b(n266), .O(n473));
  orx  g0446(.a(n473), .b(n467), .O(n474));
  orx  g0447(.a(n474), .b(n462), .O(n475));
  andx g0448(.a(n475), .b(n192), .O(n476));
  andx g0449(.a(n153), .b(n71), .O(n477));
  andx g0450(.a(n477), .b(n109), .O(n478));
  andx g0451(.a(pi12), .b(n81), .O(n479));
  andx g0452(.a(n479), .b(pi09), .O(n480));
  andx g0453(.a(n480), .b(n152), .O(n481));
  orx  g0454(.a(n481), .b(n478), .O(n482));
  andx g0455(.a(n482), .b(n29), .O(n483));
  andx g0456(.a(n266), .b(n258), .O(n484));
  andx g0457(.a(n375), .b(pi13), .O(n485));
  orx  g0458(.a(n485), .b(n484), .O(n486));
  orx  g0459(.a(n486), .b(n483), .O(n487));
  andx g0460(.a(n487), .b(n139), .O(n488));
  orx  g0461(.a(n488), .b(n476), .O(n489));
  orx  g0462(.a(n489), .b(n471), .O(n490));
  andx g0463(.a(n329), .b(n162), .O(n491));
  andx g0464(.a(n100), .b(n82), .O(n492));
  andx g0465(.a(n492), .b(n98), .O(n493));
  andx g0466(.a(n242), .b(n109), .O(n494));
  andx g0467(.a(n494), .b(n107), .O(n495));
  orx  g0468(.a(n495), .b(n493), .O(n496));
  orx  g0469(.a(n496), .b(n491), .O(n497));
  andx g0470(.a(n107), .b(n73), .O(n498));
  andx g0471(.a(n213), .b(n208), .O(n499));
  andx g0472(.a(n499), .b(n498), .O(n500));
  andx g0473(.a(n120), .b(n48), .O(n501));
  andx g0474(.a(n100), .b(n81), .O(n502));
  andx g0475(.a(n502), .b(n501), .O(n503));
  andx g0476(.a(n503), .b(n310), .O(n504));
  andx g0477(.a(n120), .b(pi05), .O(n505));
  andx g0478(.a(n505), .b(n314), .O(n506));
  andx g0479(.a(n506), .b(n502), .O(n507));
  orx  g0480(.a(n507), .b(n504), .O(n508));
  orx  g0481(.a(n508), .b(n500), .O(n509));
  orx  g0482(.a(n509), .b(n497), .O(n510));
  andx g0483(.a(n385), .b(n41), .O(n511));
  andx g0484(.a(n511), .b(n95), .O(n512));
  orx  g0485(.a(n512), .b(n387), .O(n513));
  andx g0486(.a(n513), .b(n452), .O(n514));
  andx g0487(.a(n103), .b(n28), .O(n515));
  orx  g0488(.a(n515), .b(n492), .O(n516));
  andx g0489(.a(n516), .b(n260), .O(n517));
  orx  g0490(.a(n517), .b(n514), .O(n518));
  andx g0491(.a(n515), .b(n98), .O(n519));
  andx g0492(.a(n283), .b(n109), .O(n520));
  andx g0493(.a(n520), .b(n107), .O(n521));
  orx  g0494(.a(n521), .b(n519), .O(n522));
  orx  g0495(.a(n298), .b(n79), .O(n523));
  andx g0496(.a(n523), .b(n188), .O(n524));
  orx  g0497(.a(n524), .b(n522), .O(n525));
  orx  g0498(.a(n525), .b(n518), .O(n526));
  orx  g0499(.a(n526), .b(n510), .O(n527));
  andx g0500(.a(n163), .b(n71), .O(n528));
  andx g0501(.a(n528), .b(n30), .O(n529));
  orx  g0502(.a(n529), .b(n172), .O(n530));
  andx g0503(.a(n530), .b(n126), .O(n531));
  andx g0504(.a(n230), .b(n35), .O(n532));
  andx g0505(.a(pi10), .b(n28), .O(n533));
  andx g0506(.a(n533), .b(pi08), .O(n534));
  andx g0507(.a(n33), .b(n532), .O(n535));
  andx g0508(.a(n532), .b(n123), .O(n536));
  orx  g0509(.a(n536), .b(n535), .O(n537));
  orx  g0510(.a(n537), .b(n531), .O(n538));
  andx g0511(.a(n344), .b(n126), .O(n539));
  andx g0512(.a(n539), .b(n36), .O(n540));
  andx g0513(.a(n529), .b(n126), .O(n541));
  andx g0514(.a(n541), .b(n36), .O(n542));
  orx  g0515(.a(n542), .b(n540), .O(n543));
  orx  g0516(.a(n543), .b(n538), .O(n544));
  orx  g0517(.a(n473), .b(n333), .O(n545));
  andx g0518(.a(n545), .b(n323), .O(n546));
  andx g0519(.a(n311), .b(n302), .O(n547));
  andx g0520(.a(n310), .b(pi13), .O(n548));
  andx g0521(.a(n548), .b(n547), .O(n549));
  andx g0522(.a(n315), .b(n302), .O(n550));
  andx g0523(.a(n314), .b(pi13), .O(n551));
  andx g0524(.a(n551), .b(n550), .O(n552));
  orx  g0525(.a(n552), .b(n549), .O(n553));
  orx  g0526(.a(n529), .b(n33), .O(n554));
  andx g0527(.a(n554), .b(n175), .O(n555));
  orx  g0528(.a(n555), .b(n553), .O(n556));
  orx  g0529(.a(n556), .b(n546), .O(n557));
  orx  g0530(.a(n557), .b(n544), .O(n558));
  orx  g0531(.a(n558), .b(n527), .O(n559));
  orx  g0532(.a(n559), .b(n490), .O(n560));
  orx  g0533(.a(n560), .b(n459), .O(n561));
  orx  g0534(.a(n561), .b(n250), .O(po00));
  invx g0535(.a(pi01), .O(n563));
  andx g0536(.a(pi02), .b(n563), .O(n564));
  andx g0537(.a(n564), .b(pi00), .O(n565));
  andx g0538(.a(n190), .b(pi03), .O(n566));
  andx g0539(.a(n566), .b(n565), .O(n567));
  andx g0540(.a(n567), .b(n464), .O(n568));
  andx g0541(.a(n253), .b(pi00), .O(n569));
  orx  g0542(.a(pi05), .b(n37), .O(n570));
  andx g0543(.a(n570), .b(n569), .O(n571));
  andx g0544(.a(n571), .b(n69), .O(n572));
  orx  g0545(.a(n572), .b(n568), .O(n573));
  andx g0546(.a(n569), .b(n38), .O(n574));
  andx g0547(.a(n574), .b(n203), .O(n575));
  andx g0548(.a(n565), .b(n30), .O(n576));
  andx g0549(.a(n576), .b(n383), .O(n577));
  orx  g0550(.a(n577), .b(n575), .O(n578));
  orx  g0551(.a(n578), .b(n573), .O(n579));
  andx g0552(.a(pi05), .b(n563), .O(n580));
  andx g0553(.a(n580), .b(pi02), .O(n581));
  andx g0554(.a(n581), .b(pi13), .O(n582));
  andx g0555(.a(pi09), .b(pi08), .O(n583));
  invx g0556(.a(n583), .O(n584));
  andx g0557(.a(n110), .b(pi07), .O(n585));
  andx g0558(.a(n585), .b(n584), .O(n586));
  andx g0559(.a(n586), .b(n582), .O(n587));
  andx g0560(.a(pi03), .b(pi02), .O(n588));
  andx g0561(.a(n588), .b(pi00), .O(n589));
  andx g0562(.a(n41), .b(pi04), .O(n590));
  andx g0563(.a(n590), .b(n563), .O(n591));
  andx g0564(.a(n591), .b(n589), .O(n592));
  andx g0565(.a(n592), .b(n460), .O(n593));
  orx  g0566(.a(n593), .b(n587), .O(n594));
  andx g0567(.a(n230), .b(n178), .O(n595));
  andx g0568(.a(n100), .b(pi11), .O(n596));
  andx g0569(.a(n596), .b(n420), .O(n597));
  andx g0570(.a(n597), .b(n595), .O(n598));
  orx  g0571(.a(n598), .b(n373), .O(n599));
  orx  g0572(.a(n599), .b(n594), .O(n600));
  orx  g0573(.a(n600), .b(n579), .O(n601));
  orx  g0574(.a(n418), .b(n127), .O(n602));
  andx g0575(.a(n203), .b(n44), .O(n603));
  orx  g0576(.a(n603), .b(n384), .O(n604));
  orx  g0577(.a(n604), .b(n602), .O(n605));
  andx g0578(.a(n123), .b(n44), .O(n606));
  andx g0579(.a(pi05), .b(pi03), .O(n607));
  andx g0580(.a(n607), .b(n36), .O(n608));
  andx g0581(.a(n608), .b(n298), .O(n609));
  orx  g0582(.a(n609), .b(n606), .O(n610));
  orx  g0583(.a(n338), .b(n54), .O(n611));
  orx  g0584(.a(n611), .b(n610), .O(n612));
  orx  g0585(.a(n612), .b(n605), .O(n613));
  orx  g0586(.a(n613), .b(n601), .O(n614));
  andx g0587(.a(n188), .b(pi13), .O(n615));
  andx g0588(.a(n615), .b(n547), .O(n616));
  orx  g0589(.a(n616), .b(n539), .O(n617));
  orx  g0590(.a(n617), .b(n306), .O(n618));
  andx g0591(.a(n597), .b(n581), .O(n619));
  andx g0592(.a(n588), .b(pi01), .O(n620));
  andx g0593(.a(pi07), .b(pi05), .O(n621));
  andx g0594(.a(n621), .b(n37), .O(n622));
  andx g0595(.a(n622), .b(n620), .O(n623));
  andx g0596(.a(n623), .b(n104), .O(n624));
  orx  g0597(.a(n624), .b(n619), .O(n625));
  andx g0598(.a(n571), .b(n280), .O(n626));
  andx g0599(.a(n608), .b(n422), .O(n627));
  orx  g0600(.a(n627), .b(n626), .O(n628));
  orx  g0601(.a(n628), .b(n625), .O(n629));
  orx  g0602(.a(n629), .b(n618), .O(n630));
  andx g0603(.a(n44), .b(n33), .O(n631));
  andx g0604(.a(n567), .b(n460), .O(n632));
  orx  g0605(.a(n632), .b(n631), .O(n633));
  orx  g0606(.a(n633), .b(n537), .O(n634));
  andx g0607(.a(n277), .b(n34), .O(n635));
  andx g0608(.a(n173), .b(n153), .O(n636));
  andx g0609(.a(n636), .b(n82), .O(n637));
  andx g0610(.a(n637), .b(n635), .O(n638));
  orx  g0611(.a(n638), .b(n541), .O(n639));
  andx g0612(.a(n592), .b(n467), .O(n640));
  orx  g0613(.a(n640), .b(n377), .O(n641));
  orx  g0614(.a(n641), .b(n639), .O(n642));
  orx  g0615(.a(n642), .b(n634), .O(n643));
  orx  g0616(.a(n643), .b(n630), .O(n644));
  orx  g0617(.a(n644), .b(n614), .O(n645));
  andx g0618(.a(n167), .b(n49), .O(n646));
  andx g0619(.a(n297), .b(n264), .O(n647));
  orx  g0620(.a(n647), .b(n87), .O(n648));
  andx g0621(.a(n648), .b(n646), .O(n649));
  orx  g0622(.a(n503), .b(n413), .O(n650));
  orx  g0623(.a(n650), .b(n402), .O(n651));
  andx g0624(.a(n651), .b(n188), .O(n652));
  orx  g0625(.a(n652), .b(n649), .O(n653));
  orx  g0626(.a(n653), .b(n92), .O(n654));
  andx g0627(.a(n100), .b(n83), .O(n655));
  orx  g0628(.a(n655), .b(n102), .O(n656));
  andx g0629(.a(n533), .b(pi07), .O(n657));
  andx g0630(.a(n657), .b(n596), .O(n658));
  orx  g0631(.a(n658), .b(n656), .O(n659));
  andx g0632(.a(n659), .b(n595), .O(n660));
  orx  g0633(.a(n660), .b(n118), .O(n661));
  orx  g0634(.a(n467), .b(n335), .O(n662));
  andx g0635(.a(n662), .b(n567), .O(n663));
  andx g0636(.a(n141), .b(pi04), .O(n664));
  andx g0637(.a(n664), .b(n146), .O(n665));
  andx g0638(.a(n664), .b(n143), .O(n666));
  orx  g0639(.a(n666), .b(n665), .O(n667));
  andx g0640(.a(n151), .b(pi04), .O(n668));
  andx g0641(.a(n668), .b(n154), .O(n669));
  andx g0642(.a(n147), .b(pi04), .O(n670));
  andx g0643(.a(n670), .b(n146), .O(n671));
  orx  g0644(.a(n671), .b(n669), .O(n672));
  orx  g0645(.a(n672), .b(n667), .O(n673));
  andx g0646(.a(n673), .b(n635), .O(n674));
  orx  g0647(.a(n674), .b(n663), .O(n675));
  orx  g0648(.a(n675), .b(n661), .O(n676));
  orx  g0649(.a(n676), .b(n654), .O(n677));
  orx  g0650(.a(n677), .b(n645), .O(n678));
  andx g0651(.a(n668), .b(n480), .O(n679));
  orx  g0652(.a(n477), .b(n234), .O(n680));
  andx g0653(.a(n108), .b(pi04), .O(n681));
  andx g0654(.a(n681), .b(n680), .O(n682));
  andx g0655(.a(n180), .b(pi04), .O(n683));
  andx g0656(.a(n683), .b(n362), .O(n684));
  andx g0657(.a(n255), .b(pi04), .O(n685));
  andx g0658(.a(n685), .b(n272), .O(n686));
  orx  g0659(.a(n686), .b(n684), .O(n687));
  orx  g0660(.a(n687), .b(n682), .O(n688));
  orx  g0661(.a(n688), .b(n679), .O(n689));
  andx g0662(.a(n689), .b(n635), .O(n690));
  orx  g0663(.a(n348), .b(n312), .O(n691));
  andx g0664(.a(n691), .b(n188), .O(n692));
  andx g0665(.a(n646), .b(n80), .O(n693));
  orx  g0666(.a(n693), .b(n692), .O(n694));
  andx g0667(.a(n685), .b(n266), .O(n695));
  orx  g0668(.a(n695), .b(n224), .O(n696));
  andx g0669(.a(n696), .b(n635), .O(n697));
  orx  g0670(.a(n697), .b(n496), .O(n698));
  orx  g0671(.a(n698), .b(n694), .O(n699));
  orx  g0672(.a(n699), .b(n690), .O(n700));
  andx g0673(.a(n569), .b(n29), .O(n701));
  andx g0674(.a(n570), .b(n108), .O(n702));
  andx g0675(.a(n702), .b(n680), .O(n703));
  andx g0676(.a(n151), .b(n37), .O(n704));
  andx g0677(.a(n704), .b(n480), .O(n705));
  andx g0678(.a(n570), .b(n255), .O(n706));
  andx g0679(.a(n706), .b(n272), .O(n707));
  andx g0680(.a(n362), .b(n209), .O(n708));
  orx  g0681(.a(n708), .b(n707), .O(n709));
  orx  g0682(.a(n709), .b(n705), .O(n710));
  orx  g0683(.a(n710), .b(n703), .O(n711));
  andx g0684(.a(n711), .b(n701), .O(n712));
  andx g0685(.a(n592), .b(n193), .O(n713));
  orx  g0686(.a(n592), .b(n567), .O(n714));
  andx g0687(.a(n714), .b(n162), .O(n715));
  orx  g0688(.a(n715), .b(n713), .O(n716));
  andx g0689(.a(n716), .b(n328), .O(n717));
  orx  g0690(.a(n717), .b(n712), .O(n718));
  orx  g0691(.a(n718), .b(n700), .O(n719));
  orx  g0692(.a(n172), .b(n164), .O(n720));
  andx g0693(.a(n720), .b(n44), .O(n721));
  orx  g0694(.a(n576), .b(n228), .O(n722));
  andx g0695(.a(n171), .b(n28), .O(n723));
  andx g0696(.a(n723), .b(n230), .O(n724));
  andx g0697(.a(n724), .b(n722), .O(n725));
  orx  g0698(.a(n725), .b(n721), .O(n726));
  orx  g0699(.a(n473), .b(n195), .O(n727));
  andx g0700(.a(n727), .b(n567), .O(n728));
  andx g0701(.a(n592), .b(n335), .O(n729));
  orx  g0702(.a(n729), .b(n728), .O(n730));
  orx  g0703(.a(n730), .b(n726), .O(n731));
  andx g0704(.a(n714), .b(n280), .O(n732));
  andx g0705(.a(n608), .b(n87), .O(n733));
  orx  g0706(.a(n733), .b(n732), .O(n734));
  andx g0707(.a(n714), .b(n461), .O(n735));
  andx g0708(.a(n439), .b(n52), .O(n736));
  andx g0709(.a(n622), .b(n146), .O(n737));
  orx  g0710(.a(n737), .b(n736), .O(n738));
  andx g0711(.a(n563), .b(pi00), .O(n739));
  andx g0712(.a(n739), .b(n29), .O(n740));
  andx g0713(.a(n740), .b(pi02), .O(n741));
  andx g0714(.a(n741), .b(n738), .O(n742));
  orx  g0715(.a(n742), .b(n735), .O(n743));
  orx  g0716(.a(n743), .b(n734), .O(n744));
  orx  g0717(.a(n744), .b(n731), .O(n745));
  orx  g0718(.a(pi11), .b(n81), .O(n746));
  andx g0719(.a(n327), .b(n746), .O(n747));
  orx  g0720(.a(n99), .b(n28), .O(n748));
  andx g0721(.a(n748), .b(n32), .O(n749));
  orx  g0722(.a(n749), .b(n747), .O(n750));
  andx g0723(.a(n750), .b(n230), .O(n751));
  andx g0724(.a(n751), .b(n576), .O(n752));
  andx g0725(.a(n714), .b(n69), .O(n753));
  orx  g0726(.a(n753), .b(n752), .O(n754));
  andx g0727(.a(n141), .b(pi05), .O(n755));
  andx g0728(.a(n755), .b(n143), .O(n756));
  andx g0729(.a(n756), .b(n701), .O(n757));
  andx g0730(.a(n141), .b(n37), .O(n758));
  andx g0731(.a(n758), .b(n569), .O(n759));
  andx g0732(.a(n759), .b(n279), .O(n760));
  orx  g0733(.a(n760), .b(n757), .O(n761));
  andx g0734(.a(n49), .b(pi02), .O(n762));
  andx g0735(.a(n550), .b(n29), .O(n763));
  andx g0736(.a(n763), .b(n762), .O(n764));
  orx  g0737(.a(n764), .b(n761), .O(n765));
  orx  g0738(.a(n765), .b(n754), .O(n766));
  andx g0739(.a(n135), .b(n132), .O(n767));
  orx  g0740(.a(n767), .b(n442), .O(n768));
  orx  g0741(.a(n768), .b(n522), .O(n769));
  andx g0742(.a(n77), .b(pi05), .O(n770));
  andx g0743(.a(n770), .b(n37), .O(n771));
  andx g0744(.a(n771), .b(n620), .O(n772));
  orx  g0745(.a(n772), .b(n215), .O(n773));
  orx  g0746(.a(n452), .b(n217), .O(n774));
  andx g0747(.a(n774), .b(n773), .O(n775));
  orx  g0748(.a(n775), .b(n500), .O(n776));
  orx  g0749(.a(n776), .b(n769), .O(n777));
  orx  g0750(.a(n777), .b(n766), .O(n778));
  orx  g0751(.a(n778), .b(n745), .O(n779));
  andx g0752(.a(n574), .b(n530), .O(n780));
  andx g0753(.a(n259), .b(n104), .O(n781));
  andx g0754(.a(n515), .b(n259), .O(n782));
  orx  g0755(.a(n782), .b(n781), .O(n783));
  orx  g0756(.a(n783), .b(n780), .O(n784));
  andx g0757(.a(n727), .b(n592), .O(n785));
  andx g0758(.a(n151), .b(pi05), .O(n786));
  andx g0759(.a(n786), .b(n154), .O(n787));
  andx g0760(.a(n147), .b(pi05), .O(n788));
  andx g0761(.a(n788), .b(n146), .O(n789));
  orx  g0762(.a(n789), .b(n787), .O(n790));
  andx g0763(.a(n790), .b(n701), .O(n791));
  orx  g0764(.a(n791), .b(n785), .O(n792));
  orx  g0765(.a(n792), .b(n784), .O(n793));
  andx g0766(.a(n229), .b(n153), .O(n794));
  andx g0767(.a(n794), .b(n82), .O(n795));
  andx g0768(.a(n795), .b(n701), .O(n796));
  andx g0769(.a(n786), .b(n480), .O(n797));
  andx g0770(.a(n797), .b(n701), .O(n798));
  orx  g0771(.a(n798), .b(n796), .O(n799));
  andx g0772(.a(n259), .b(n102), .O(n800));
  andx g0773(.a(n623), .b(n515), .O(n801));
  orx  g0774(.a(n801), .b(n800), .O(n802));
  orx  g0775(.a(n802), .b(n799), .O(n803));
  andx g0776(.a(n143), .b(n29), .O(n804));
  andx g0777(.a(n804), .b(n759), .O(n805));
  andx g0778(.a(n574), .b(n164), .O(n806));
  orx  g0779(.a(n806), .b(n805), .O(n807));
  andx g0780(.a(n100), .b(n78), .O(n808));
  andx g0781(.a(n808), .b(n581), .O(n809));
  andx g0782(.a(n755), .b(n146), .O(n810));
  andx g0783(.a(n810), .b(n701), .O(n811));
  orx  g0784(.a(n811), .b(n809), .O(n812));
  orx  g0785(.a(n812), .b(n807), .O(n813));
  orx  g0786(.a(n813), .b(n803), .O(n814));
  orx  g0787(.a(n814), .b(n793), .O(n815));
  andx g0788(.a(n714), .b(n407), .O(n816));
  andx g0789(.a(n103), .b(n72), .O(n817));
  orx  g0790(.a(n817), .b(n808), .O(n818));
  andx g0791(.a(n818), .b(n595), .O(n819));
  orx  g0792(.a(n819), .b(n816), .O(n820));
  andx g0793(.a(n656), .b(n581), .O(n821));
  orx  g0794(.a(n339), .b(n202), .O(n822));
  andx g0795(.a(n822), .b(n230), .O(n823));
  andx g0796(.a(n823), .b(n576), .O(n824));
  orx  g0797(.a(n824), .b(n821), .O(n825));
  orx  g0798(.a(n825), .b(n820), .O(n826));
  andx g0799(.a(n620), .b(n242), .O(n827));
  andx g0800(.a(n620), .b(n114), .O(n828));
  orx  g0801(.a(n828), .b(n827), .O(n829));
  andx g0802(.a(n622), .b(pi13), .O(n830));
  andx g0803(.a(n830), .b(n829), .O(n831));
  andx g0804(.a(n512), .b(n452), .O(n832));
  andx g0805(.a(n492), .b(n259), .O(n833));
  orx  g0806(.a(n833), .b(n832), .O(n834));
  orx  g0807(.a(n834), .b(n831), .O(n835));
  andx g0808(.a(n99), .b(pi09), .O(n836));
  andx g0809(.a(n836), .b(pi07), .O(n837));
  andx g0810(.a(n837), .b(n230), .O(n838));
  orx  g0811(.a(n838), .b(n441), .O(n839));
  andx g0812(.a(n839), .b(n576), .O(n840));
  andx g0813(.a(n608), .b(n80), .O(n841));
  orx  g0814(.a(n841), .b(n840), .O(n842));
  orx  g0815(.a(n842), .b(n835), .O(n843));
  orx  g0816(.a(n843), .b(n826), .O(n844));
  orx  g0817(.a(n844), .b(n815), .O(n845));
  orx  g0818(.a(n845), .b(n779), .O(n846));
  orx  g0819(.a(n846), .b(n719), .O(n847));
  orx  g0820(.a(n847), .b(n678), .O(po01));
  andx g0821(.a(n705), .b(n701), .O(n849));
  andx g0822(.a(n382), .b(n240), .O(n850));
  andx g0823(.a(n850), .b(n576), .O(n851));
  orx  g0824(.a(n851), .b(n849), .O(n852));
  andx g0825(.a(n138), .b(pi00), .O(n853));
  andx g0826(.a(n853), .b(n29), .O(n854));
  andx g0827(.a(n854), .b(n481), .O(n855));
  andx g0828(.a(n153), .b(n81), .O(n856));
  andx g0829(.a(n856), .b(n466), .O(n857));
  andx g0830(.a(n590), .b(pi01), .O(n858));
  andx g0831(.a(n858), .b(n29), .O(n859));
  andx g0832(.a(n859), .b(n857), .O(n860));
  orx  g0833(.a(n860), .b(n855), .O(n861));
  orx  g0834(.a(n861), .b(n852), .O(n862));
  andx g0835(.a(n481), .b(n47), .O(n863));
  andx g0836(.a(n145), .b(n81), .O(n864));
  andx g0837(.a(n864), .b(n466), .O(n865));
  andx g0838(.a(n865), .b(n859), .O(n866));
  orx  g0839(.a(n866), .b(n863), .O(n867));
  andx g0840(.a(n110), .b(pi09), .O(n868));
  andx g0841(.a(n868), .b(n350), .O(n869));
  andx g0842(.a(n869), .b(n551), .O(n870));
  andx g0843(.a(n49), .b(n36), .O(n871));
  andx g0844(.a(n74), .b(n81), .O(n872));
  andx g0845(.a(n872), .b(n466), .O(n873));
  andx g0846(.a(n873), .b(n871), .O(n874));
  orx  g0847(.a(n874), .b(n870), .O(n875));
  orx  g0848(.a(n875), .b(n867), .O(n876));
  orx  g0849(.a(n876), .b(n862), .O(n877));
  andx g0850(.a(pi10), .b(pi09), .O(n878));
  andx g0851(.a(n878), .b(pi08), .O(n879));
  andx g0852(.a(n879), .b(n209), .O(n880));
  andx g0853(.a(n880), .b(n57), .O(n881));
  andx g0854(.a(n879), .b(n361), .O(n882));
  andx g0855(.a(n882), .b(n35), .O(n883));
  orx  g0856(.a(n883), .b(n881), .O(n884));
  andx g0857(.a(n884), .b(n30), .O(n885));
  orx  g0858(.a(n858), .b(n323), .O(n886));
  andx g0859(.a(n886), .b(n856), .O(n887));
  andx g0860(.a(n871), .b(n868), .O(n888));
  orx  g0861(.a(n888), .b(n887), .O(n889));
  andx g0862(.a(n406), .b(n29), .O(n890));
  andx g0863(.a(n890), .b(n889), .O(n891));
  orx  g0864(.a(n891), .b(n885), .O(n892));
  orx  g0865(.a(n892), .b(n877), .O(n893));
  andx g0866(.a(n381), .b(pi08), .O(n894));
  andx g0867(.a(n894), .b(n209), .O(n895));
  andx g0868(.a(n569), .b(n30), .O(n896));
  andx g0869(.a(n896), .b(n895), .O(n897));
  andx g0870(.a(n865), .b(n278), .O(n898));
  orx  g0871(.a(n898), .b(n897), .O(n899));
  andx g0872(.a(n502), .b(n466), .O(n900));
  andx g0873(.a(n900), .b(n139), .O(n901));
  andx g0874(.a(n569), .b(n181), .O(n902));
  andx g0875(.a(n894), .b(n30), .O(n903));
  andx g0876(.a(n903), .b(n902), .O(n904));
  orx  g0877(.a(n904), .b(n901), .O(n905));
  orx  g0878(.a(n905), .b(n899), .O(n906));
  andx g0879(.a(n59), .b(pi01), .O(n907));
  andx g0880(.a(n907), .b(n277), .O(n908));
  andx g0881(.a(n908), .b(pi12), .O(n909));
  andx g0882(.a(n99), .b(n81), .O(n910));
  andx g0883(.a(n910), .b(pi09), .O(n911));
  andx g0884(.a(n911), .b(n240), .O(n912));
  andx g0885(.a(n912), .b(n909), .O(n913));
  andx g0886(.a(n438), .b(pi02), .O(n914));
  andx g0887(.a(n327), .b(pi07), .O(n915));
  andx g0888(.a(n915), .b(n103), .O(n916));
  andx g0889(.a(n916), .b(n914), .O(n917));
  orx  g0890(.a(n917), .b(n913), .O(n918));
  andx g0891(.a(n655), .b(n581), .O(n919));
  andx g0892(.a(n49), .b(pi00), .O(n920));
  andx g0893(.a(n920), .b(n30), .O(n921));
  andx g0894(.a(n921), .b(n895), .O(n922));
  orx  g0895(.a(n922), .b(n919), .O(n923));
  orx  g0896(.a(n923), .b(n918), .O(n924));
  orx  g0897(.a(n924), .b(n906), .O(n925));
  andx g0898(.a(n868), .b(n347), .O(n926));
  andx g0899(.a(n926), .b(n107), .O(n927));
  andx g0900(.a(n909), .b(n895), .O(n928));
  orx  g0901(.a(n928), .b(n927), .O(n929));
  andx g0902(.a(n574), .b(n529), .O(n930));
  andx g0903(.a(n879), .b(n180), .O(n931));
  andx g0904(.a(n858), .b(n30), .O(n932));
  andx g0905(.a(n932), .b(n931), .O(n933));
  orx  g0906(.a(n933), .b(n930), .O(n934));
  orx  g0907(.a(n934), .b(n929), .O(n935));
  andx g0908(.a(n900), .b(n254), .O(n936));
  andx g0909(.a(n503), .b(n95), .O(n937));
  orx  g0910(.a(n937), .b(n936), .O(n938));
  andx g0911(.a(n37), .b(pi02), .O(n939));
  andx g0912(.a(n939), .b(n563), .O(n940));
  andx g0913(.a(n940), .b(pi13), .O(n941));
  andx g0914(.a(n72), .b(pi06), .O(n942));
  andx g0915(.a(n942), .b(n868), .O(n943));
  andx g0916(.a(n943), .b(n941), .O(n944));
  orx  g0917(.a(pi06), .b(n41), .O(n945));
  andx g0918(.a(n945), .b(n72), .O(n946));
  andx g0919(.a(n946), .b(n139), .O(n947));
  andx g0920(.a(n103), .b(pi09), .O(n948));
  andx g0921(.a(n948), .b(n947), .O(n949));
  orx  g0922(.a(n949), .b(n944), .O(n950));
  orx  g0923(.a(n950), .b(n938), .O(n951));
  orx  g0924(.a(n951), .b(n935), .O(n952));
  orx  g0925(.a(n952), .b(n925), .O(n953));
  orx  g0926(.a(n953), .b(n893), .O(n954));
  andx g0927(.a(n382), .b(n109), .O(n955));
  andx g0928(.a(n853), .b(n30), .O(n956));
  andx g0929(.a(n63), .b(pi00), .O(n957));
  andx g0930(.a(n957), .b(n30), .O(n958));
  orx  g0931(.a(n958), .b(n956), .O(n959));
  andx g0932(.a(n959), .b(n955), .O(n960));
  andx g0933(.a(n177), .b(pi00), .O(n961));
  andx g0934(.a(n961), .b(n681), .O(n962));
  andx g0935(.a(n569), .b(n240), .O(n963));
  orx  g0936(.a(n963), .b(n962), .O(n964));
  andx g0937(.a(n964), .b(n164), .O(n965));
  orx  g0938(.a(n965), .b(n960), .O(n966));
  andx g0939(.a(n911), .b(n109), .O(n967));
  andx g0940(.a(n967), .b(n959), .O(n968));
  andx g0941(.a(n921), .b(n912), .O(n969));
  andx g0942(.a(n119), .b(n82), .O(n970));
  andx g0943(.a(n970), .b(n962), .O(n971));
  orx  g0944(.a(n971), .b(n969), .O(n972));
  orx  g0945(.a(n972), .b(n968), .O(n973));
  andx g0946(.a(n569), .b(n358), .O(n974));
  andx g0947(.a(n974), .b(n164), .O(n975));
  andx g0948(.a(n921), .b(n850), .O(n976));
  andx g0949(.a(n702), .b(n569), .O(n977));
  andx g0950(.a(n977), .b(n970), .O(n978));
  orx  g0951(.a(n978), .b(n976), .O(n979));
  orx  g0952(.a(n979), .b(n975), .O(n980));
  orx  g0953(.a(n980), .b(n973), .O(n981));
  orx  g0954(.a(n981), .b(n966), .O(n982));
  andx g0955(.a(n311), .b(n107), .O(n983));
  andx g0956(.a(n406), .b(n179), .O(n984));
  orx  g0957(.a(n984), .b(n983), .O(n985));
  andx g0958(.a(n985), .b(n868), .O(n986));
  andx g0959(.a(n882), .b(n853), .O(n987));
  andx g0960(.a(n920), .b(n880), .O(n988));
  orx  g0961(.a(n988), .b(n987), .O(n989));
  andx g0962(.a(n989), .b(n193), .O(n990));
  orx  g0963(.a(n990), .b(n986), .O(n991));
  andx g0964(.a(n879), .b(n193), .O(n992));
  andx g0965(.a(n571), .b(n180), .O(n993));
  andx g0966(.a(n961), .b(n683), .O(n994));
  andx g0967(.a(n957), .b(n361), .O(n995));
  orx  g0968(.a(n995), .b(n994), .O(n996));
  orx  g0969(.a(n996), .b(n993), .O(n997));
  andx g0970(.a(n997), .b(n992), .O(n998));
  andx g0971(.a(n501), .b(n266), .O(n999));
  orx  g0972(.a(n999), .b(n465), .O(n1000));
  andx g0973(.a(n1000), .b(n323), .O(n1001));
  orx  g0974(.a(n1001), .b(n998), .O(n1002));
  orx  g0975(.a(n1002), .b(n991), .O(n1003));
  orx  g0976(.a(n1003), .b(n982), .O(n1004));
  orx  g0977(.a(n1004), .b(n954), .O(n1005));
  andx g0978(.a(n74), .b(pi10), .O(n1006));
  orx  g0979(.a(pi05), .b(pi04), .O(n1007));
  orx  g0980(.a(n48), .b(n41), .O(n1008));
  andx g0981(.a(n1008), .b(pi02), .O(n1009));
  andx g0982(.a(n1009), .b(n1007), .O(n1010));
  orx  g0983(.a(n1010), .b(n168), .O(n1011));
  andx g0984(.a(n1011), .b(n1006), .O(n1012));
  andx g0985(.a(n582), .b(n110), .O(n1013));
  orx  g0986(.a(n1013), .b(n1012), .O(n1014));
  andx g0987(.a(n583), .b(n77), .O(n1015));
  orx  g0988(.a(n1015), .b(n915), .O(n1016));
  andx g0989(.a(n1016), .b(n1014), .O(n1017));
  andx g0990(.a(n931), .b(n73), .O(n1018));
  andx g0991(.a(n1018), .b(n287), .O(n1019));
  andx g0992(.a(n920), .b(n29), .O(n1020));
  andx g0993(.a(n51), .b(pi09), .O(n1021));
  andx g0994(.a(n1021), .b(n256), .O(n1022));
  orx  g0995(.a(n1022), .b(n787), .O(n1023));
  andx g0996(.a(n1023), .b(n1020), .O(n1024));
  orx  g0997(.a(n1024), .b(n1019), .O(n1025));
  orx  g0998(.a(n1020), .b(n701), .O(n1026));
  andx g0999(.a(n1026), .b(n797), .O(n1027));
  andx g1000(.a(n1018), .b(n941), .O(n1028));
  orx  g1001(.a(n1028), .b(n1027), .O(n1029));
  orx  g1002(.a(n1029), .b(n1025), .O(n1030));
  orx  g1003(.a(n1030), .b(n1017), .O(n1031));
  andx g1004(.a(n879), .b(n119), .O(n1032));
  orx  g1005(.a(n996), .b(n989), .O(n1033));
  andx g1006(.a(n1033), .b(n1032), .O(n1034));
  andx g1007(.a(n607), .b(pi01), .O(n1035));
  andx g1008(.a(n1035), .b(pi13), .O(n1036));
  orx  g1009(.a(n1036), .b(n548), .O(n1037));
  andx g1010(.a(n1037), .b(n311), .O(n1038));
  andx g1011(.a(n551), .b(n315), .O(n1039));
  andx g1012(.a(n858), .b(pi13), .O(n1040));
  andx g1013(.a(n1040), .b(n406), .O(n1041));
  orx  g1014(.a(n1041), .b(n1039), .O(n1042));
  orx  g1015(.a(n1042), .b(n1038), .O(n1043));
  andx g1016(.a(n1043), .b(n868), .O(n1044));
  orx  g1017(.a(n1044), .b(n1034), .O(n1045));
  orx  g1018(.a(n1045), .b(n1031), .O(n1046));
  andx g1019(.a(n1021), .b(n258), .O(n1047));
  orx  g1020(.a(n1047), .b(n155), .O(n1048));
  andx g1021(.a(n1048), .b(n47), .O(n1049));
  andx g1022(.a(n909), .b(n850), .O(n1050));
  andx g1023(.a(n912), .b(n576), .O(n1051));
  orx  g1024(.a(n1051), .b(n1050), .O(n1052));
  orx  g1025(.a(n1052), .b(n1049), .O(n1053));
  orx  g1026(.a(n909), .b(n576), .O(n1054));
  andx g1027(.a(n1054), .b(n880), .O(n1055));
  andx g1028(.a(n957), .b(n29), .O(n1056));
  orx  g1029(.a(n1056), .b(n854), .O(n1057));
  andx g1030(.a(n1057), .b(n1047), .O(n1058));
  orx  g1031(.a(n1058), .b(n1055), .O(n1059));
  orx  g1032(.a(n1059), .b(n1053), .O(n1060));
  andx g1033(.a(n967), .b(n228), .O(n1061));
  andx g1034(.a(n57), .b(n30), .O(n1062));
  andx g1035(.a(n1062), .b(n912), .O(n1063));
  orx  g1036(.a(n1063), .b(n1061), .O(n1064));
  andx g1037(.a(n961), .b(n29), .O(n1065));
  andx g1038(.a(n1021), .b(n685), .O(n1066));
  orx  g1039(.a(n1066), .b(n669), .O(n1067));
  andx g1040(.a(n1067), .b(n1065), .O(n1068));
  orx  g1041(.a(n1068), .b(n1064), .O(n1069));
  orx  g1042(.a(n608), .b(n188), .O(n1070));
  orx  g1043(.a(n1070), .b(n1010), .O(n1071));
  andx g1044(.a(n1071), .b(n84), .O(n1072));
  orx  g1045(.a(n1062), .b(n576), .O(n1073));
  andx g1046(.a(n1073), .b(n895), .O(n1074));
  orx  g1047(.a(n1074), .b(n1072), .O(n1075));
  orx  g1048(.a(n1075), .b(n1069), .O(n1076));
  orx  g1049(.a(n1076), .b(n1060), .O(n1077));
  andx g1050(.a(n871), .b(n29), .O(n1078));
  orx  g1051(.a(n1078), .b(n1040), .O(n1079));
  andx g1052(.a(n1079), .b(n943), .O(n1080));
  andx g1053(.a(n894), .b(n361), .O(n1081));
  andx g1054(.a(n1081), .b(n959), .O(n1082));
  orx  g1055(.a(n1082), .b(n1080), .O(n1083));
  orx  g1056(.a(n797), .b(n787), .O(n1084));
  orx  g1057(.a(n908), .b(n741), .O(n1085));
  andx g1058(.a(n1085), .b(n1084), .O(n1086));
  orx  g1059(.a(n1086), .b(n508), .O(n1087));
  orx  g1060(.a(n1087), .b(n1083), .O(n1088));
  andx g1061(.a(n1037), .b(n926), .O(n1089));
  andx g1062(.a(n1065), .b(n679), .O(n1090));
  andx g1063(.a(n1056), .b(n481), .O(n1091));
  orx  g1064(.a(n1091), .b(n1090), .O(n1092));
  orx  g1065(.a(n1092), .b(n1089), .O(n1093));
  andx g1066(.a(n945), .b(n201), .O(n1094));
  andx g1067(.a(n1094), .b(n239), .O(n1095));
  andx g1068(.a(n1095), .b(n868), .O(n1096));
  orx  g1069(.a(n287), .b(n179), .O(n1097));
  andx g1070(.a(n1097), .b(n943), .O(n1098));
  orx  g1071(.a(n1098), .b(n1096), .O(n1099));
  orx  g1072(.a(n1099), .b(n1093), .O(n1100));
  orx  g1073(.a(n1100), .b(n1088), .O(n1101));
  orx  g1074(.a(n1101), .b(n1077), .O(n1102));
  andx g1075(.a(n57), .b(n29), .O(n1103));
  andx g1076(.a(n1103), .b(n787), .O(n1104));
  andx g1077(.a(n406), .b(n323), .O(n1105));
  andx g1078(.a(n266), .b(n163), .O(n1106));
  andx g1079(.a(n1106), .b(n1105), .O(n1107));
  orx  g1080(.a(n1107), .b(n1104), .O(n1108));
  andx g1081(.a(n96), .b(pi09), .O(n1109));
  andx g1082(.a(n1109), .b(n139), .O(n1110));
  andx g1083(.a(n1110), .b(n502), .O(n1111));
  andx g1084(.a(n1035), .b(n503), .O(n1112));
  orx  g1085(.a(n1112), .b(n1111), .O(n1113));
  orx  g1086(.a(n1113), .b(n1108), .O(n1114));
  andx g1087(.a(n1022), .b(n908), .O(n1115));
  orx  g1088(.a(n1115), .b(n200), .O(n1116));
  andx g1089(.a(n857), .b(n278), .O(n1117));
  andx g1090(.a(n836), .b(n266), .O(n1118));
  andx g1091(.a(n1118), .b(n1105), .O(n1119));
  orx  g1092(.a(n1119), .b(n1117), .O(n1120));
  orx  g1093(.a(n1120), .b(n1116), .O(n1121));
  orx  g1094(.a(n1121), .b(n1114), .O(n1122));
  andx g1095(.a(n1022), .b(n701), .O(n1123));
  andx g1096(.a(n994), .b(n903), .O(n1124));
  orx  g1097(.a(n1124), .b(n1123), .O(n1125));
  andx g1098(.a(n1081), .b(n228), .O(n1126));
  andx g1099(.a(n1022), .b(n741), .O(n1127));
  orx  g1100(.a(n1127), .b(n1126), .O(n1128));
  orx  g1101(.a(n1128), .b(n1125), .O(n1129));
  andx g1102(.a(n858), .b(n464), .O(n1130));
  andx g1103(.a(n858), .b(n463), .O(n1131));
  orx  g1104(.a(n1131), .b(n1130), .O(n1132));
  andx g1105(.a(n940), .b(n900), .O(n1133));
  andx g1106(.a(n1015), .b(n1006), .O(n1134));
  andx g1107(.a(n1134), .b(n608), .O(n1135));
  orx  g1108(.a(n1135), .b(n1133), .O(n1136));
  orx  g1109(.a(n1136), .b(n1132), .O(n1137));
  orx  g1110(.a(n1137), .b(n1129), .O(n1138));
  orx  g1111(.a(n1138), .b(n1122), .O(n1139));
  andx g1112(.a(n1062), .b(n850), .O(n1140));
  andx g1113(.a(n955), .b(n228), .O(n1141));
  orx  g1114(.a(n1141), .b(n1140), .O(n1142));
  andx g1115(.a(n1057), .b(n155), .O(n1143));
  orx  g1116(.a(n1143), .b(n1142), .O(n1144));
  andx g1117(.a(n255), .b(n37), .O(n1145));
  andx g1118(.a(n1145), .b(n1021), .O(n1146));
  orx  g1119(.a(n1146), .b(n787), .O(n1147));
  andx g1120(.a(n1147), .b(n701), .O(n1148));
  andx g1121(.a(n1015), .b(n103), .O(n1149));
  orx  g1122(.a(n1149), .b(n655), .O(n1150));
  andx g1123(.a(n1150), .b(n914), .O(n1151));
  orx  g1124(.a(n1151), .b(n1148), .O(n1152));
  orx  g1125(.a(n1152), .b(n1144), .O(n1153));
  orx  g1126(.a(n1022), .b(n797), .O(n1154));
  andx g1127(.a(n1154), .b(n1103), .O(n1155));
  andx g1128(.a(n900), .b(n178), .O(n1156));
  andx g1129(.a(n1006), .b(n915), .O(n1157));
  andx g1130(.a(n1157), .b(n608), .O(n1158));
  orx  g1131(.a(n1158), .b(n1156), .O(n1159));
  orx  g1132(.a(n1159), .b(n1155), .O(n1160));
  orx  g1133(.a(n999), .b(n900), .O(n1161));
  andx g1134(.a(n1161), .b(n858), .O(n1162));
  andx g1135(.a(n1032), .b(n993), .O(n1163));
  orx  g1136(.a(n1163), .b(n1162), .O(n1164));
  orx  g1137(.a(n1164), .b(n1160), .O(n1165));
  orx  g1138(.a(n1165), .b(n1153), .O(n1166));
  orx  g1139(.a(n1166), .b(n1139), .O(n1167));
  orx  g1140(.a(n1167), .b(n1102), .O(n1168));
  orx  g1141(.a(n1168), .b(n1046), .O(n1169));
  orx  g1142(.a(n1169), .b(n1005), .O(po02));
  andx g1143(.a(n406), .b(n302), .O(n1171));
  andx g1144(.a(n1171), .b(n1040), .O(n1172));
  andx g1145(.a(n301), .b(pi10), .O(n1173));
  andx g1146(.a(n1173), .b(n401), .O(n1174));
  andx g1147(.a(n1174), .b(n548), .O(n1175));
  orx  g1148(.a(n1175), .b(n1172), .O(n1176));
  andx g1149(.a(n381), .b(n100), .O(n1177));
  andx g1150(.a(n1177), .b(n1110), .O(n1178));
  andx g1151(.a(pi11), .b(pi10), .O(n1179));
  andx g1152(.a(n1179), .b(n100), .O(n1180));
  andx g1153(.a(n1180), .b(n399), .O(n1181));
  orx  g1154(.a(n1181), .b(n1178), .O(n1182));
  orx  g1155(.a(n1182), .b(n1176), .O(n1183));
  andx g1156(.a(n301), .b(n81), .O(n1184));
  andx g1157(.a(n1184), .b(n501), .O(n1185));
  andx g1158(.a(n1185), .b(n107), .O(n1186));
  andx g1159(.a(n1177), .b(n506), .O(n1187));
  orx  g1160(.a(n1187), .b(n1186), .O(n1188));
  andx g1161(.a(n1171), .b(n941), .O(n1189));
  andx g1162(.a(n1020), .b(n795), .O(n1190));
  orx  g1163(.a(n1190), .b(n1189), .O(n1191));
  orx  g1164(.a(n1191), .b(n1188), .O(n1192));
  orx  g1165(.a(n1192), .b(n1183), .O(n1193));
  andx g1166(.a(n153), .b(pi10), .O(n1194));
  andx g1167(.a(n1194), .b(n256), .O(n1195));
  andx g1168(.a(n1195), .b(n1020), .O(n1196));
  andx g1169(.a(n71), .b(n77), .O(n1197));
  andx g1170(.a(n1197), .b(pi06), .O(n1198));
  andx g1171(.a(n1198), .b(n154), .O(n1199));
  andx g1172(.a(n1199), .b(n859), .O(n1200));
  orx  g1173(.a(n1200), .b(n1196), .O(n1201));
  andx g1174(.a(n1171), .b(n287), .O(n1202));
  andx g1175(.a(n1173), .b(n915), .O(n1203));
  andx g1176(.a(n1203), .b(n582), .O(n1204));
  orx  g1177(.a(n1204), .b(n1202), .O(n1205));
  orx  g1178(.a(n1205), .b(n1201), .O(n1206));
  andx g1179(.a(n1065), .b(n686), .O(n1207));
  andx g1180(.a(n1056), .b(n294), .O(n1208));
  orx  g1181(.a(n1208), .b(n1207), .O(n1209));
  andx g1182(.a(n1145), .b(n272), .O(n1210));
  andx g1183(.a(n1210), .b(n701), .O(n1211));
  orx  g1184(.a(n1211), .b(n806), .O(n1212));
  orx  g1185(.a(n1212), .b(n1209), .O(n1213));
  orx  g1186(.a(n1213), .b(n1206), .O(n1214));
  orx  g1187(.a(n1214), .b(n1193), .O(n1215));
  andx g1188(.a(n854), .b(n294), .O(n1216));
  andx g1189(.a(n914), .b(n658), .O(n1217));
  orx  g1190(.a(n1217), .b(n1216), .O(n1218));
  andx g1191(.a(n1184), .b(n466), .O(n1219));
  andx g1192(.a(n1219), .b(n1078), .O(n1220));
  orx  g1193(.a(n1220), .b(n796), .O(n1221));
  orx  g1194(.a(n1221), .b(n1218), .O(n1222));
  andx g1195(.a(n397), .b(pi06), .O(n1223));
  andx g1196(.a(n1223), .b(n1173), .O(n1224));
  andx g1197(.a(n1224), .b(n1078), .O(n1225));
  andx g1198(.a(n583), .b(n193), .O(n1226));
  andx g1199(.a(n1226), .b(n994), .O(n1227));
  orx  g1200(.a(n1227), .b(n1225), .O(n1228));
  andx g1201(.a(n1065), .b(n637), .O(n1229));
  orx  g1202(.a(n1229), .b(n367), .O(n1230));
  orx  g1203(.a(n1230), .b(n1228), .O(n1231));
  orx  g1204(.a(n1231), .b(n1222), .O(n1232));
  andx g1205(.a(n130), .b(n71), .O(n1233));
  andx g1206(.a(n1233), .b(n30), .O(n1234));
  andx g1207(.a(n1234), .b(n977), .O(n1235));
  andx g1208(.a(n272), .b(n256), .O(n1236));
  andx g1209(.a(n1236), .b(n701), .O(n1237));
  orx  g1210(.a(n1237), .b(n1235), .O(n1238));
  andx g1211(.a(n945), .b(n397), .O(n1239));
  andx g1212(.a(n1239), .b(n1173), .O(n1240));
  andx g1213(.a(n1240), .b(n239), .O(n1241));
  andx g1214(.a(n657), .b(n421), .O(n1242));
  orx  g1215(.a(n608), .b(n168), .O(n1243));
  andx g1216(.a(n1243), .b(n1242), .O(n1244));
  orx  g1217(.a(n1244), .b(n1241), .O(n1245));
  orx  g1218(.a(n1245), .b(n1238), .O(n1246));
  andx g1219(.a(n1242), .b(n1010), .O(n1247));
  orx  g1220(.a(n1247), .b(n619), .O(n1248));
  andx g1221(.a(n1173), .b(n406), .O(n1249));
  andx g1222(.a(n1249), .b(n941), .O(n1250));
  andx g1223(.a(n421), .b(n83), .O(n1251));
  andx g1224(.a(n1251), .b(n608), .O(n1252));
  orx  g1225(.a(n1252), .b(n1250), .O(n1253));
  orx  g1226(.a(n1253), .b(n1248), .O(n1254));
  orx  g1227(.a(n1254), .b(n1246), .O(n1255));
  orx  g1228(.a(n1255), .b(n1232), .O(n1256));
  orx  g1229(.a(n1256), .b(n1215), .O(n1257));
  orx  g1230(.a(n1097), .b(n940), .O(n1258));
  andx g1231(.a(n163), .b(n103), .O(n1259));
  andx g1232(.a(n1259), .b(n942), .O(n1260));
  andx g1233(.a(n1260), .b(n1258), .O(n1261));
  andx g1234(.a(n163), .b(pi08), .O(n1262));
  andx g1235(.a(n1262), .b(n209), .O(n1263));
  andx g1236(.a(n1233), .b(n240), .O(n1264));
  orx  g1237(.a(n1264), .b(n1263), .O(n1265));
  andx g1238(.a(n528), .b(n209), .O(n1266));
  orx  g1239(.a(n1266), .b(n1265), .O(n1267));
  andx g1240(.a(n1267), .b(n1062), .O(n1268));
  orx  g1241(.a(n1268), .b(n1261), .O(n1269));
  andx g1242(.a(n1173), .b(n311), .O(n1270));
  andx g1243(.a(n1179), .b(pi09), .O(n1271));
  andx g1244(.a(n1271), .b(n347), .O(n1272));
  andx g1245(.a(n1272), .b(n73), .O(n1273));
  orx  g1246(.a(n1273), .b(n1270), .O(n1274));
  andx g1247(.a(n1274), .b(n548), .O(n1275));
  andx g1248(.a(n1173), .b(n1042), .O(n1276));
  orx  g1249(.a(n1276), .b(n1275), .O(n1277));
  orx  g1250(.a(n1277), .b(n1269), .O(n1278));
  andx g1251(.a(n1267), .b(n1054), .O(n1279));
  andx g1252(.a(n528), .b(n361), .O(n1280));
  andx g1253(.a(n1233), .b(n109), .O(n1281));
  orx  g1254(.a(n1281), .b(n1280), .O(n1282));
  andx g1255(.a(n1262), .b(n361), .O(n1283));
  orx  g1256(.a(n1283), .b(n1282), .O(n1284));
  andx g1257(.a(n1284), .b(n228), .O(n1285));
  orx  g1258(.a(n1285), .b(n1279), .O(n1286));
  orx  g1259(.a(n48), .b(n37), .O(n1287));
  andx g1260(.a(n621), .b(n1287), .O(n1288));
  andx g1261(.a(n1035), .b(n72), .O(n1289));
  andx g1262(.a(n1289), .b(n1288), .O(n1290));
  orx  g1263(.a(n1290), .b(n947), .O(n1291));
  andx g1264(.a(n1291), .b(n1259), .O(n1292));
  andx g1265(.a(n942), .b(n272), .O(n1293));
  andx g1266(.a(n1194), .b(n472), .O(n1294));
  andx g1267(.a(n406), .b(n154), .O(n1295));
  orx  g1268(.a(n1295), .b(n1294), .O(n1296));
  orx  g1269(.a(n1296), .b(n1293), .O(n1297));
  andx g1270(.a(n1297), .b(n278), .O(n1298));
  orx  g1271(.a(n1298), .b(n1292), .O(n1299));
  orx  g1272(.a(n1299), .b(n1286), .O(n1300));
  orx  g1273(.a(n1300), .b(n1278), .O(n1301));
  orx  g1274(.a(n1301), .b(n1257), .O(n1302));
  andx g1275(.a(n1224), .b(n1097), .O(n1303));
  orx  g1276(.a(n1236), .b(n1195), .O(n1304));
  andx g1277(.a(n1304), .b(n1103), .O(n1305));
  orx  g1278(.a(n1305), .b(n1303), .O(n1306));
  andx g1279(.a(n1185), .b(n1037), .O(n1307));
  orx  g1280(.a(n608), .b(n199), .O(n1308));
  andx g1281(.a(n29), .b(pi05), .O(n1309));
  andx g1282(.a(n1309), .b(n1308), .O(n1310));
  andx g1283(.a(n1310), .b(n1203), .O(n1311));
  orx  g1284(.a(n1311), .b(n1307), .O(n1312));
  orx  g1285(.a(n1312), .b(n1306), .O(n1313));
  andx g1286(.a(n1282), .b(n959), .O(n1314));
  andx g1287(.a(n1304), .b(n1085), .O(n1315));
  orx  g1288(.a(n1315), .b(n1314), .O(n1316));
  andx g1289(.a(n1095), .b(n302), .O(n1317));
  orx  g1290(.a(n1317), .b(n553), .O(n1318));
  orx  g1291(.a(n1318), .b(n1316), .O(n1319));
  orx  g1292(.a(n1319), .b(n1313), .O(n1320));
  andx g1293(.a(n1194), .b(n258), .O(n1321));
  andx g1294(.a(n1321), .b(n1057), .O(n1322));
  orx  g1295(.a(n1321), .b(n294), .O(n1323));
  andx g1296(.a(n1323), .b(n47), .O(n1324));
  andx g1297(.a(n1219), .b(n1097), .O(n1325));
  orx  g1298(.a(n1325), .b(n1324), .O(n1326));
  orx  g1299(.a(n1326), .b(n1322), .O(n1327));
  andx g1300(.a(n1179), .b(n28), .O(n1328));
  andx g1301(.a(n1328), .b(n755), .O(n1329));
  andx g1302(.a(n1329), .b(n1073), .O(n1330));
  andx g1303(.a(n590), .b(pi02), .O(n1331));
  orx  g1304(.a(n1331), .b(n188), .O(n1332));
  andx g1305(.a(n1332), .b(n29), .O(n1333));
  andx g1306(.a(n1333), .b(n1203), .O(n1334));
  orx  g1307(.a(n1334), .b(n1330), .O(n1335));
  orx  g1308(.a(n1224), .b(n1219), .O(n1336));
  andx g1309(.a(n1336), .b(n941), .O(n1337));
  orx  g1310(.a(n1103), .b(n741), .O(n1338));
  andx g1311(.a(n1338), .b(n795), .O(n1339));
  orx  g1312(.a(n1339), .b(n1337), .O(n1340));
  orx  g1313(.a(n1340), .b(n1335), .O(n1341));
  orx  g1314(.a(n1341), .b(n1327), .O(n1342));
  orx  g1315(.a(n1342), .b(n1320), .O(n1343));
  andx g1316(.a(n193), .b(n68), .O(n1344));
  orx  g1317(.a(n1344), .b(n195), .O(n1345));
  andx g1318(.a(n1345), .b(n858), .O(n1346));
  orx  g1319(.a(n921), .b(n896), .O(n1347));
  andx g1320(.a(n1347), .b(n1266), .O(n1348));
  orx  g1321(.a(n1348), .b(n1346), .O(n1349));
  andx g1322(.a(n871), .b(n74), .O(n1350));
  andx g1323(.a(n858), .b(n100), .O(n1351));
  orx  g1324(.a(n1351), .b(n1350), .O(n1352));
  andx g1325(.a(n1271), .b(n942), .O(n1353));
  andx g1326(.a(n1353), .b(n1352), .O(n1354));
  orx  g1327(.a(n1035), .b(n95), .O(n1355));
  andx g1328(.a(n1355), .b(pi13), .O(n1356));
  andx g1329(.a(n1356), .b(n1174), .O(n1357));
  orx  g1330(.a(n1357), .b(n1354), .O(n1358));
  orx  g1331(.a(n1358), .b(n1349), .O(n1359));
  andx g1332(.a(n1270), .b(n1036), .O(n1360));
  andx g1333(.a(n1249), .b(n287), .O(n1361));
  orx  g1334(.a(n1361), .b(n1360), .O(n1362));
  andx g1335(.a(n1199), .b(n278), .O(n1363));
  andx g1336(.a(n1295), .b(n859), .O(n1364));
  orx  g1337(.a(n1364), .b(n1363), .O(n1365));
  orx  g1338(.a(n1365), .b(n1362), .O(n1366));
  andx g1339(.a(n1272), .b(n498), .O(n1367));
  andx g1340(.a(n1356), .b(n547), .O(n1368));
  orx  g1341(.a(n1368), .b(n1367), .O(n1369));
  orx  g1342(.a(n1369), .b(n1366), .O(n1370));
  orx  g1343(.a(n1370), .b(n1359), .O(n1371));
  andx g1344(.a(n1328), .b(n142), .O(n1372));
  orx  g1345(.a(n1372), .b(n1283), .O(n1373));
  andx g1346(.a(n1373), .b(n959), .O(n1374));
  orx  g1347(.a(n1329), .b(n1263), .O(n1375));
  andx g1348(.a(n1375), .b(n896), .O(n1376));
  orx  g1349(.a(n1376), .b(n1374), .O(n1377));
  andx g1350(.a(n1173), .b(n1095), .O(n1378));
  andx g1351(.a(n1265), .b(n921), .O(n1379));
  orx  g1352(.a(n1379), .b(n1378), .O(n1380));
  orx  g1353(.a(n1380), .b(n1377), .O(n1381));
  andx g1354(.a(n1251), .b(n1011), .O(n1382));
  orx  g1355(.a(n854), .b(n47), .O(n1383));
  andx g1356(.a(n1383), .b(n273), .O(n1384));
  orx  g1357(.a(n1384), .b(n1382), .O(n1385));
  orx  g1358(.a(n1331), .b(n199), .O(n1386));
  orx  g1359(.a(n1386), .b(n1070), .O(n1387));
  andx g1360(.a(n421), .b(n78), .O(n1388));
  andx g1361(.a(n1388), .b(n1387), .O(n1389));
  orx  g1362(.a(n994), .b(n902), .O(n1390));
  andx g1363(.a(n1390), .b(n529), .O(n1391));
  orx  g1364(.a(n1391), .b(n1389), .O(n1392));
  orx  g1365(.a(n1392), .b(n1385), .O(n1393));
  orx  g1366(.a(n1393), .b(n1381), .O(n1394));
  orx  g1367(.a(n1394), .b(n1371), .O(n1395));
  andx g1368(.a(n1293), .b(n859), .O(n1396));
  andx g1369(.a(n1194), .b(n706), .O(n1397));
  andx g1370(.a(n1397), .b(n701), .O(n1398));
  orx  g1371(.a(n1398), .b(n1396), .O(n1399));
  andx g1372(.a(n1194), .b(n685), .O(n1400));
  andx g1373(.a(n1400), .b(n1065), .O(n1401));
  andx g1374(.a(n1056), .b(n273), .O(n1402));
  orx  g1375(.a(n1402), .b(n1401), .O(n1403));
  orx  g1376(.a(n1403), .b(n1399), .O(n1404));
  andx g1377(.a(n914), .b(n550), .O(n1405));
  andx g1378(.a(n1249), .b(n1078), .O(n1406));
  orx  g1379(.a(n1406), .b(n1405), .O(n1407));
  andx g1380(.a(n1386), .b(n422), .O(n1408));
  andx g1381(.a(n1294), .b(n859), .O(n1409));
  orx  g1382(.a(n1409), .b(n1408), .O(n1410));
  orx  g1383(.a(n1410), .b(n1407), .O(n1411));
  orx  g1384(.a(n1411), .b(n1404), .O(n1412));
  andx g1385(.a(n1219), .b(n1040), .O(n1413));
  andx g1386(.a(n596), .b(n83), .O(n1414));
  andx g1387(.a(n1414), .b(n914), .O(n1415));
  orx  g1388(.a(n1415), .b(n1413), .O(n1416));
  andx g1389(.a(n1328), .b(n30), .O(n1417));
  andx g1390(.a(n1417), .b(n759), .O(n1418));
  andx g1391(.a(n1344), .b(n323), .O(n1419));
  orx  g1392(.a(n1419), .b(n1418), .O(n1420));
  orx  g1393(.a(n1420), .b(n1416), .O(n1421));
  andx g1394(.a(n1236), .b(n1020), .O(n1422));
  andx g1395(.a(n1224), .b(n1040), .O(n1423));
  orx  g1396(.a(n1423), .b(n1422), .O(n1424));
  andx g1397(.a(n460), .b(n323), .O(n1425));
  andx g1398(.a(n1219), .b(n239), .O(n1426));
  orx  g1399(.a(n1426), .b(n1425), .O(n1427));
  orx  g1400(.a(n1427), .b(n1424), .O(n1428));
  orx  g1401(.a(n1428), .b(n1421), .O(n1429));
  orx  g1402(.a(n1429), .b(n1412), .O(n1430));
  andx g1403(.a(n961), .b(n664), .O(n1431));
  andx g1404(.a(n1431), .b(n1417), .O(n1432));
  andx g1405(.a(n1329), .b(n909), .O(n1433));
  orx  g1406(.a(n1433), .b(n1432), .O(n1434));
  andx g1407(.a(n1226), .b(n902), .O(n1435));
  andx g1408(.a(n1372), .b(n228), .O(n1436));
  orx  g1409(.a(n1436), .b(n1435), .O(n1437));
  orx  g1410(.a(n1437), .b(n1434), .O(n1438));
  andx g1411(.a(n908), .b(n795), .O(n1439));
  andx g1412(.a(n1329), .b(n921), .O(n1440));
  orx  g1413(.a(n1440), .b(n1439), .O(n1441));
  andx g1414(.a(n1249), .b(n179), .O(n1442));
  andx g1415(.a(n1234), .b(n962), .O(n1443));
  orx  g1416(.a(n1443), .b(n1442), .O(n1444));
  orx  g1417(.a(n1444), .b(n1441), .O(n1445));
  orx  g1418(.a(n1445), .b(n1438), .O(n1446));
  andx g1419(.a(n1171), .b(n1078), .O(n1447));
  andx g1420(.a(n858), .b(n460), .O(n1448));
  orx  g1421(.a(n1448), .b(n1447), .O(n1449));
  andx g1422(.a(n1414), .b(n581), .O(n1450));
  andx g1423(.a(n1070), .b(n422), .O(n1451));
  orx  g1424(.a(n1451), .b(n1450), .O(n1452));
  orx  g1425(.a(n1452), .b(n1449), .O(n1453));
  orx  g1426(.a(n657), .b(n78), .O(n1454));
  andx g1427(.a(n596), .b(n581), .O(n1455));
  andx g1428(.a(n1455), .b(n1454), .O(n1456));
  andx g1429(.a(n1171), .b(n179), .O(n1457));
  orx  g1430(.a(n1457), .b(n1456), .O(n1458));
  orx  g1431(.a(n915), .b(n201), .O(n1459));
  andx g1432(.a(n1173), .b(n914), .O(n1460));
  andx g1433(.a(n1460), .b(n1459), .O(n1461));
  andx g1434(.a(n1270), .b(n107), .O(n1462));
  orx  g1435(.a(n1462), .b(n1461), .O(n1463));
  orx  g1436(.a(n1463), .b(n1458), .O(n1464));
  orx  g1437(.a(n1464), .b(n1453), .O(n1465));
  orx  g1438(.a(n1465), .b(n1446), .O(n1466));
  orx  g1439(.a(n1466), .b(n1430), .O(n1467));
  orx  g1440(.a(n1467), .b(n1395), .O(n1468));
  orx  g1441(.a(n1468), .b(n1343), .O(n1469));
  orx  g1442(.a(n1469), .b(n1302), .O(po03));
  andx g1443(.a(n89), .b(n36), .O(n1471));
  andx g1444(.a(n138), .b(pi02), .O(n1472));
  orx  g1445(.a(n1472), .b(n1471), .O(n1473));
  andx g1446(.a(n872), .b(n505), .O(n1474));
  andx g1447(.a(n1474), .b(n1473), .O(n1475));
  andx g1448(.a(n139), .b(n103), .O(n1476));
  andx g1449(.a(n1476), .b(n303), .O(n1477));
  orx  g1450(.a(n1477), .b(n1475), .O(n1478));
  andx g1451(.a(n438), .b(pi03), .O(n1479));
  andx g1452(.a(n1479), .b(n440), .O(n1480));
  andx g1453(.a(n30), .b(n563), .O(n1481));
  andx g1454(.a(n36), .b(pi00), .O(n1482));
  andx g1455(.a(n1482), .b(n1481), .O(n1483));
  andx g1456(.a(n1483), .b(n1480), .O(n1484));
  andx g1457(.a(n1471), .b(n647), .O(n1485));
  orx  g1458(.a(n1485), .b(n1484), .O(n1486));
  orx  g1459(.a(n1486), .b(n1478), .O(n1487));
  andx g1460(.a(n96), .b(n71), .O(n1488));
  orx  g1461(.a(n1488), .b(n1223), .O(n1489));
  andx g1462(.a(n1489), .b(n1476), .O(n1490));
  andx g1463(.a(n63), .b(n563), .O(n1491));
  andx g1464(.a(n1491), .b(n428), .O(n1492));
  orx  g1465(.a(n1492), .b(n1490), .O(n1493));
  andx g1466(.a(n397), .b(n41), .O(n1494));
  andx g1467(.a(n1494), .b(n1476), .O(n1495));
  orx  g1468(.a(n1495), .b(n1111), .O(n1496));
  orx  g1469(.a(n1496), .b(n1493), .O(n1497));
  orx  g1470(.a(n1497), .b(n1487), .O(n1498));
  andx g1471(.a(n229), .b(pi03), .O(n1499));
  orx  g1472(.a(n837), .b(n122), .O(n1500));
  andx g1473(.a(n1500), .b(n576), .O(n1501));
  andx g1474(.a(n1483), .b(n747), .O(n1502));
  orx  g1475(.a(n1502), .b(n1501), .O(n1503));
  andx g1476(.a(n1503), .b(n1499), .O(n1504));
  orx  g1477(.a(n908), .b(n278), .O(n1505));
  andx g1478(.a(n477), .b(n240), .O(n1506));
  orx  g1479(.a(n1236), .b(n708), .O(n1507));
  orx  g1480(.a(n1507), .b(n1506), .O(n1508));
  andx g1481(.a(n1508), .b(n1505), .O(n1509));
  orx  g1482(.a(n1509), .b(n1504), .O(n1510));
  orx  g1483(.a(n1510), .b(n1498), .O(n1511));
  andx g1484(.a(n229), .b(n59), .O(n1512));
  andx g1485(.a(n1512), .b(n202), .O(n1513));
  andx g1486(.a(n1513), .b(n1062), .O(n1514));
  orx  g1487(.a(n1514), .b(n495), .O(n1515));
  andx g1488(.a(n1499), .b(n202), .O(n1516));
  andx g1489(.a(n1516), .b(n1483), .O(n1517));
  andx g1490(.a(n229), .b(pi04), .O(n1518));
  andx g1491(.a(n1518), .b(n254), .O(n1519));
  andx g1492(.a(n1519), .b(n597), .O(n1520));
  orx  g1493(.a(n1520), .b(n1517), .O(n1521));
  orx  g1494(.a(n1521), .b(n1515), .O(n1522));
  andx g1495(.a(n961), .b(n30), .O(n1523));
  andx g1496(.a(n1518), .b(n202), .O(n1524));
  andx g1497(.a(n1524), .b(n1523), .O(n1525));
  andx g1498(.a(n1480), .b(n576), .O(n1526));
  orx  g1499(.a(n1526), .b(n1525), .O(n1527));
  andx g1500(.a(n1491), .b(pi13), .O(n1528));
  andx g1501(.a(n1528), .b(n550), .O(n1529));
  andx g1502(.a(n1499), .b(n382), .O(n1530));
  andx g1503(.a(n1530), .b(n576), .O(n1531));
  orx  g1504(.a(n1531), .b(n1529), .O(n1532));
  orx  g1505(.a(n1532), .b(n1527), .O(n1533));
  orx  g1506(.a(n1533), .b(n1522), .O(n1534));
  andx g1507(.a(n494), .b(n287), .O(n1535));
  orx  g1508(.a(n1535), .b(n800), .O(n1536));
  andx g1509(.a(n907), .b(n276), .O(n1537));
  orx  g1510(.a(n1537), .b(n323), .O(n1538));
  andx g1511(.a(n1538), .b(n267), .O(n1539));
  andx g1512(.a(n1472), .b(n647), .O(n1540));
  orx  g1513(.a(n1540), .b(n1539), .O(n1541));
  orx  g1514(.a(n1541), .b(n1536), .O(n1542));
  andx g1515(.a(n1516), .b(n576), .O(n1543));
  andx g1516(.a(n1499), .b(n339), .O(n1544));
  andx g1517(.a(n1544), .b(n1483), .O(n1545));
  orx  g1518(.a(n1545), .b(n1543), .O(n1546));
  andx g1519(.a(n1518), .b(n382), .O(n1547));
  andx g1520(.a(n1547), .b(n1523), .O(n1548));
  andx g1521(.a(n1512), .b(n382), .O(n1549));
  andx g1522(.a(n1549), .b(n1062), .O(n1550));
  orx  g1523(.a(n1550), .b(n1548), .O(n1551));
  orx  g1524(.a(n1551), .b(n1546), .O(n1552));
  orx  g1525(.a(n1552), .b(n1542), .O(n1553));
  orx  g1526(.a(n1553), .b(n1534), .O(n1554));
  orx  g1527(.a(n1554), .b(n1511), .O(n1555));
  andx g1528(.a(n438), .b(pi04), .O(n1556));
  andx g1529(.a(n1556), .b(n440), .O(n1557));
  orx  g1530(.a(n534), .b(n528), .O(n1558));
  orx  g1531(.a(n1558), .b(n1500), .O(n1559));
  orx  g1532(.a(n28), .b(pi08), .O(n1560));
  andx g1533(.a(n1560), .b(n171), .O(n1561));
  orx  g1534(.a(n1561), .b(n339), .O(n1562));
  orx  g1535(.a(n1562), .b(n1559), .O(n1563));
  andx g1536(.a(n1563), .b(n1518), .O(n1564));
  orx  g1537(.a(n1564), .b(n1557), .O(n1565));
  andx g1538(.a(n1565), .b(n1523), .O(n1566));
  andx g1539(.a(n505), .b(n502), .O(n1567));
  andx g1540(.a(n621), .b(n584), .O(n1568));
  orx  g1541(.a(n1568), .b(n315), .O(n1569));
  andx g1542(.a(n1569), .b(n103), .O(n1570));
  orx  g1543(.a(n1570), .b(n1567), .O(n1571));
  andx g1544(.a(n1571), .b(n1491), .O(n1572));
  andx g1545(.a(n438), .b(n59), .O(n1573));
  andx g1546(.a(n1573), .b(n440), .O(n1574));
  andx g1547(.a(n1562), .b(n1512), .O(n1575));
  orx  g1548(.a(n1575), .b(n1574), .O(n1576));
  andx g1549(.a(n1576), .b(n1062), .O(n1577));
  andx g1550(.a(n1559), .b(n1512), .O(n1578));
  andx g1551(.a(n1578), .b(n1062), .O(n1579));
  orx  g1552(.a(n1579), .b(n1577), .O(n1580));
  orx  g1553(.a(n1580), .b(n1572), .O(n1581));
  orx  g1554(.a(n1581), .b(n1566), .O(n1582));
  orx  g1555(.a(n1582), .b(n1555), .O(n1583));
  andx g1556(.a(n102), .b(pi06), .O(n1584));
  orx  g1557(.a(n1584), .b(n900), .O(n1585));
  andx g1558(.a(n291), .b(n101), .O(n1586));
  orx  g1559(.a(n1586), .b(n1585), .O(n1587));
  andx g1560(.a(n1587), .b(n139), .O(n1588));
  andx g1561(.a(n566), .b(n56), .O(n1589));
  orx  g1562(.a(n818), .b(n659), .O(n1590));
  andx g1563(.a(n1590), .b(n1589), .O(n1591));
  orx  g1564(.a(n1561), .b(n1558), .O(n1592));
  andx g1565(.a(n1592), .b(n576), .O(n1593));
  orx  g1566(.a(n1561), .b(n382), .O(n1594));
  orx  g1567(.a(n1594), .b(n749), .O(n1595));
  andx g1568(.a(n1595), .b(n1483), .O(n1596));
  orx  g1569(.a(n1596), .b(n1593), .O(n1597));
  andx g1570(.a(n1597), .b(n1499), .O(n1598));
  orx  g1571(.a(n1598), .b(n1591), .O(n1599));
  orx  g1572(.a(n1599), .b(n1588), .O(n1600));
  orx  g1573(.a(n422), .b(n298), .O(n1601));
  orx  g1574(.a(n1601), .b(n88), .O(n1602));
  andx g1575(.a(n1602), .b(n1331), .O(n1603));
  orx  g1576(.a(n287), .b(n107), .O(n1604));
  andx g1577(.a(n1604), .b(n115), .O(n1605));
  andx g1578(.a(n920), .b(n268), .O(n1606));
  orx  g1579(.a(n1606), .b(n1605), .O(n1607));
  andx g1580(.a(n1589), .b(n48), .O(n1608));
  andx g1581(.a(n1608), .b(n597), .O(n1609));
  andx g1582(.a(n406), .b(n103), .O(n1610));
  andx g1583(.a(n942), .b(n103), .O(n1611));
  orx  g1584(.a(n1611), .b(n1610), .O(n1612));
  andx g1585(.a(n1612), .b(n139), .O(n1613));
  orx  g1586(.a(n1613), .b(n1609), .O(n1614));
  orx  g1587(.a(n1614), .b(n1607), .O(n1615));
  orx  g1588(.a(n1615), .b(n1603), .O(n1616));
  andx g1589(.a(n240), .b(n234), .O(n1617));
  orx  g1590(.a(n1617), .b(n1508), .O(n1618));
  andx g1591(.a(n1618), .b(n1020), .O(n1619));
  orx  g1592(.a(n810), .b(n756), .O(n1620));
  orx  g1593(.a(n1620), .b(n1617), .O(n1621));
  orx  g1594(.a(n795), .b(n789), .O(n1622));
  orx  g1595(.a(n1622), .b(n1084), .O(n1623));
  orx  g1596(.a(n1623), .b(n1621), .O(n1624));
  andx g1597(.a(n1624), .b(n1505), .O(n1625));
  orx  g1598(.a(n1625), .b(n1619), .O(n1626));
  orx  g1599(.a(n1626), .b(n1616), .O(n1627));
  andx g1600(.a(n361), .b(n208), .O(n1628));
  orx  g1601(.a(n1628), .b(n520), .O(n1629));
  andx g1602(.a(n1629), .b(n393), .O(n1630));
  orx  g1603(.a(n1630), .b(n834), .O(n1631));
  andx g1604(.a(n1479), .b(n52), .O(n1632));
  andx g1605(.a(n621), .b(pi03), .O(n1633));
  andx g1606(.a(n1633), .b(n146), .O(n1634));
  orx  g1607(.a(n1634), .b(n1632), .O(n1635));
  andx g1608(.a(n1635), .b(n740), .O(n1636));
  andx g1609(.a(n1622), .b(n1020), .O(n1637));
  orx  g1610(.a(n1637), .b(n1636), .O(n1638));
  orx  g1611(.a(n1638), .b(n1631), .O(n1639));
  andx g1612(.a(n1538), .b(n265), .O(n1640));
  orx  g1613(.a(n1640), .b(n521), .O(n1641));
  andx g1614(.a(n1499), .b(n837), .O(n1642));
  andx g1615(.a(n1642), .b(n1483), .O(n1643));
  andx g1616(.a(n1544), .b(n576), .O(n1644));
  orx  g1617(.a(n1644), .b(n1643), .O(n1645));
  orx  g1618(.a(n1645), .b(n1641), .O(n1646));
  orx  g1619(.a(n372), .b(n112), .O(n1647));
  andx g1620(.a(n1647), .b(n1604), .O(n1648));
  orx  g1621(.a(n1648), .b(n783), .O(n1649));
  orx  g1622(.a(n1649), .b(n1646), .O(n1650));
  orx  g1623(.a(n1650), .b(n1639), .O(n1651));
  andx g1624(.a(n1556), .b(n52), .O(n1652));
  andx g1625(.a(n145), .b(pi05), .O(n1653));
  andx g1626(.a(n1653), .b(n223), .O(n1654));
  orx  g1627(.a(n1654), .b(n1652), .O(n1655));
  andx g1628(.a(n1655), .b(n1065), .O(n1656));
  andx g1629(.a(n1473), .b(n763), .O(n1657));
  orx  g1630(.a(n1657), .b(n1656), .O(n1658));
  andx g1631(.a(n1084), .b(n1020), .O(n1659));
  andx g1632(.a(n1473), .b(n1006), .O(n1660));
  andx g1633(.a(n1660), .b(n1569), .O(n1661));
  orx  g1634(.a(n1661), .b(n1659), .O(n1662));
  orx  g1635(.a(n1662), .b(n1658), .O(n1663));
  andx g1636(.a(n1573), .b(n52), .O(n1664));
  andx g1637(.a(n621), .b(n59), .O(n1665));
  andx g1638(.a(n1665), .b(n146), .O(n1666));
  orx  g1639(.a(n1666), .b(n1664), .O(n1667));
  andx g1640(.a(n1667), .b(n1103), .O(n1668));
  orx  g1641(.a(n1668), .b(n1317), .O(n1669));
  andx g1642(.a(n1620), .b(n1020), .O(n1670));
  orx  g1643(.a(n1670), .b(n500), .O(n1671));
  orx  g1644(.a(n1671), .b(n1669), .O(n1672));
  orx  g1645(.a(n1672), .b(n1663), .O(n1673));
  orx  g1646(.a(n1673), .b(n1651), .O(n1674));
  orx  g1647(.a(n1674), .b(n1627), .O(n1675));
  orx  g1648(.a(n1675), .b(n1600), .O(n1676));
  orx  g1649(.a(n1676), .b(n1583), .O(po04));
  andx g1650(.a(n755), .b(n382), .O(n1678));
  andx g1651(.a(n1678), .b(n896), .O(n1679));
  orx  g1652(.a(n1679), .b(n1172), .O(n1680));
  andx g1653(.a(n1065), .b(n665), .O(n1681));
  andx g1654(.a(n362), .b(n194), .O(n1682));
  andx g1655(.a(n1682), .b(n278), .O(n1683));
  orx  g1656(.a(n1683), .b(n1681), .O(n1684));
  orx  g1657(.a(n1684), .b(n1680), .O(n1685));
  orx  g1658(.a(n1189), .b(n575), .O(n1686));
  andx g1659(.a(n1678), .b(n921), .O(n1687));
  andx g1660(.a(n908), .b(n708), .O(n1688));
  orx  g1661(.a(n1688), .b(n1687), .O(n1689));
  orx  g1662(.a(n1689), .b(n1686), .O(n1690));
  orx  g1663(.a(n1690), .b(n1685), .O(n1691));
  andx g1664(.a(n681), .b(n114), .O(n1692));
  andx g1665(.a(n286), .b(n59), .O(n1693));
  andx g1666(.a(n1693), .b(n1692), .O(n1694));
  andx g1667(.a(n1692), .b(n287), .O(n1695));
  orx  g1668(.a(n1695), .b(n1694), .O(n1696));
  andx g1669(.a(n551), .b(n375), .O(n1697));
  orx  g1670(.a(n1697), .b(n805), .O(n1698));
  orx  g1671(.a(n1698), .b(n1696), .O(n1699));
  andx g1672(.a(n836), .b(pi08), .O(n1700));
  andx g1673(.a(n1700), .b(n240), .O(n1701));
  andx g1674(.a(n1701), .b(n896), .O(n1702));
  andx g1675(.a(n51), .b(pi08), .O(n1703));
  andx g1676(.a(n1703), .b(n256), .O(n1704));
  andx g1677(.a(n1704), .b(n1020), .O(n1705));
  orx  g1678(.a(n1705), .b(n1702), .O(n1706));
  andx g1679(.a(n1472), .b(n29), .O(n1707));
  andx g1680(.a(n1707), .b(n319), .O(n1708));
  andx g1681(.a(n683), .b(n208), .O(n1709));
  andx g1682(.a(n1709), .b(n393), .O(n1710));
  orx  g1683(.a(n1710), .b(n1708), .O(n1711));
  orx  g1684(.a(n1711), .b(n1706), .O(n1712));
  orx  g1685(.a(n1712), .b(n1699), .O(n1713));
  orx  g1686(.a(n1713), .b(n1691), .O(n1714));
  andx g1687(.a(n256), .b(n208), .O(n1715));
  andx g1688(.a(n1715), .b(n896), .O(n1716));
  andx g1689(.a(n685), .b(n208), .O(n1717));
  andx g1690(.a(n1717), .b(n1523), .O(n1718));
  orx  g1691(.a(n1718), .b(n1716), .O(n1719));
  andx g1692(.a(n741), .b(n708), .O(n1720));
  andx g1693(.a(n908), .b(n810), .O(n1721));
  orx  g1694(.a(n1721), .b(n1720), .O(n1722));
  orx  g1695(.a(n1722), .b(n1719), .O(n1723));
  andx g1696(.a(n854), .b(n156), .O(n1724));
  andx g1697(.a(n1171), .b(n582), .O(n1725));
  orx  g1698(.a(n1725), .b(n1724), .O(n1726));
  andx g1699(.a(n858), .b(n333), .O(n1727));
  orx  g1700(.a(n1727), .b(n360), .O(n1728));
  orx  g1701(.a(n1728), .b(n1726), .O(n1729));
  orx  g1702(.a(n1729), .b(n1723), .O(n1730));
  andx g1703(.a(n1682), .b(n859), .O(n1731));
  andx g1704(.a(n1065), .b(n684), .O(n1732));
  orx  g1705(.a(n1732), .b(n1731), .O(n1733));
  andx g1706(.a(n1103), .b(n810), .O(n1734));
  orx  g1707(.a(n1734), .b(n1447), .O(n1735));
  orx  g1708(.a(n1735), .b(n1733), .O(n1736));
  andx g1709(.a(n1715), .b(n909), .O(n1737));
  andx g1710(.a(n1331), .b(n873), .O(n1738));
  orx  g1711(.a(n1738), .b(n1737), .O(n1739));
  andx g1712(.a(n382), .b(n142), .O(n1740));
  andx g1713(.a(n1740), .b(n228), .O(n1741));
  andx g1714(.a(n1145), .b(n208), .O(n1742));
  andx g1715(.a(n1742), .b(n896), .O(n1743));
  orx  g1716(.a(n1743), .b(n1741), .O(n1744));
  orx  g1717(.a(n1744), .b(n1739), .O(n1745));
  orx  g1718(.a(n1745), .b(n1736), .O(n1746));
  orx  g1719(.a(n1746), .b(n1730), .O(n1747));
  orx  g1720(.a(n1747), .b(n1714), .O(n1748));
  orx  g1721(.a(n284), .b(n243), .O(n1749));
  orx  g1722(.a(n415), .b(n375), .O(n1750));
  orx  g1723(.a(n1750), .b(n1749), .O(n1751));
  andx g1724(.a(n1751), .b(n1707), .O(n1752));
  andx g1725(.a(n69), .b(pi08), .O(n1753));
  orx  g1726(.a(n1753), .b(n407), .O(n1754));
  andx g1727(.a(n1754), .b(n323), .O(n1755));
  orx  g1728(.a(n1755), .b(n1752), .O(n1756));
  andx g1729(.a(n961), .b(n695), .O(n1757));
  orx  g1730(.a(n1757), .b(n572), .O(n1758));
  andx g1731(.a(n1758), .b(pi08), .O(n1759));
  orx  g1732(.a(n426), .b(n370), .O(n1760));
  orx  g1733(.a(n1760), .b(n431), .O(n1761));
  andx g1734(.a(n1761), .b(n179), .O(n1762));
  orx  g1735(.a(n1762), .b(n1759), .O(n1763));
  orx  g1736(.a(n1763), .b(n1756), .O(n1764));
  orx  g1737(.a(n1701), .b(n1678), .O(n1765));
  orx  g1738(.a(n1765), .b(n1715), .O(n1766));
  andx g1739(.a(n1766), .b(n1073), .O(n1767));
  orx  g1740(.a(n156), .b(n144), .O(n1768));
  andx g1741(.a(n1703), .b(n258), .O(n1769));
  orx  g1742(.a(n1769), .b(n363), .O(n1770));
  orx  g1743(.a(n1770), .b(n1768), .O(n1771));
  andx g1744(.a(n1771), .b(n47), .O(n1772));
  orx  g1745(.a(n1772), .b(n1767), .O(n1773));
  andx g1746(.a(n551), .b(n209), .O(n1774));
  andx g1747(.a(n181), .b(n179), .O(n1775));
  orx  g1748(.a(n1775), .b(n1774), .O(n1776));
  andx g1749(.a(n1776), .b(n217), .O(n1777));
  orx  g1750(.a(n1332), .b(n608), .O(n1778));
  orx  g1751(.a(n1778), .b(n871), .O(n1779));
  andx g1752(.a(n1006), .b(n406), .O(n1780));
  andx g1753(.a(n1780), .b(n1779), .O(n1781));
  orx  g1754(.a(n1781), .b(n1777), .O(n1782));
  orx  g1755(.a(n1782), .b(n1773), .O(n1783));
  orx  g1756(.a(n1783), .b(n1764), .O(n1784));
  orx  g1757(.a(n1784), .b(n1748), .O(n1785));
  andx g1758(.a(n286), .b(n173), .O(n1786));
  andx g1759(.a(n1786), .b(n77), .O(n1787));
  orx  g1760(.a(n1787), .b(n1776), .O(n1788));
  andx g1761(.a(n1788), .b(n182), .O(n1789));
  andx g1762(.a(n1223), .b(n103), .O(n1790));
  orx  g1763(.a(n1790), .b(n1612), .O(n1791));
  orx  g1764(.a(n1791), .b(n1585), .O(n1792));
  andx g1765(.a(n570), .b(n564), .O(n1793));
  andx g1766(.a(n1793), .b(n1792), .O(n1794));
  orx  g1767(.a(n1794), .b(n1789), .O(n1795));
  orx  g1768(.a(n1790), .b(n473), .O(n1796));
  orx  g1769(.a(n1796), .b(n1585), .O(n1797));
  andx g1770(.a(n1797), .b(n858), .O(n1798));
  orx  g1771(.a(n1754), .b(n1612), .O(n1799));
  andx g1772(.a(n1799), .b(n858), .O(n1800));
  orx  g1773(.a(n1800), .b(n1798), .O(n1801));
  orx  g1774(.a(n1801), .b(n1795), .O(n1802));
  andx g1775(.a(n1769), .b(n1057), .O(n1803));
  orx  g1776(.a(n1803), .b(n1670), .O(n1804));
  andx g1777(.a(n1765), .b(n909), .O(n1805));
  orx  g1778(.a(n1070), .b(n871), .O(n1806));
  andx g1779(.a(n1006), .b(n942), .O(n1807));
  andx g1780(.a(n1807), .b(n1806), .O(n1808));
  orx  g1781(.a(n1808), .b(n1805), .O(n1809));
  orx  g1782(.a(n1809), .b(n1804), .O(n1810));
  andx g1783(.a(pi08), .b(pi07), .O(n1811));
  andx g1784(.a(n1811), .b(n48), .O(n1812));
  andx g1785(.a(n1812), .b(n272), .O(n1813));
  andx g1786(.a(n1811), .b(pi06), .O(n1814));
  andx g1787(.a(n1814), .b(n234), .O(n1815));
  orx  g1788(.a(n1815), .b(n1813), .O(n1816));
  andx g1789(.a(n1816), .b(n278), .O(n1817));
  andx g1790(.a(n1693), .b(n73), .O(n1818));
  andx g1791(.a(n1818), .b(n1709), .O(n1819));
  orx  g1792(.a(n1819), .b(n1817), .O(n1820));
  andx g1793(.a(n1026), .b(n708), .O(n1821));
  orx  g1794(.a(n1821), .b(n546), .O(n1822));
  orx  g1795(.a(n1822), .b(n1820), .O(n1823));
  orx  g1796(.a(n1823), .b(n1810), .O(n1824));
  andx g1797(.a(n920), .b(n240), .O(n1825));
  orx  g1798(.a(n1825), .b(n962), .O(n1826));
  andx g1799(.a(n1700), .b(n30), .O(n1827));
  andx g1800(.a(n1827), .b(n1826), .O(n1828));
  andx g1801(.a(n1057), .b(n363), .O(n1829));
  andx g1802(.a(n1171), .b(n29), .O(n1830));
  andx g1803(.a(n1830), .b(n1778), .O(n1831));
  orx  g1804(.a(n1831), .b(n1829), .O(n1832));
  orx  g1805(.a(n1832), .b(n1828), .O(n1833));
  andx g1806(.a(n1223), .b(n1006), .O(n1834));
  andx g1807(.a(n29), .b(pi06), .O(n1835));
  andx g1808(.a(n1835), .b(n113), .O(n1836));
  andx g1809(.a(n1836), .b(n67), .O(n1837));
  orx  g1810(.a(n1837), .b(n1834), .O(n1838));
  andx g1811(.a(n1838), .b(n1806), .O(n1839));
  andx g1812(.a(n258), .b(n208), .O(n1840));
  andx g1813(.a(n1840), .b(n959), .O(n1841));
  orx  g1814(.a(n1841), .b(n1839), .O(n1842));
  orx  g1815(.a(n655), .b(n586), .O(n1843));
  andx g1816(.a(n1843), .b(n1786), .O(n1844));
  orx  g1817(.a(n1704), .b(n756), .O(n1845));
  andx g1818(.a(n1845), .b(n1338), .O(n1846));
  orx  g1819(.a(n1846), .b(n1844), .O(n1847));
  orx  g1820(.a(n1847), .b(n1842), .O(n1848));
  orx  g1821(.a(n1848), .b(n1833), .O(n1849));
  orx  g1822(.a(n1849), .b(n1824), .O(n1850));
  andx g1823(.a(n1806), .b(n873), .O(n1851));
  orx  g1824(.a(n1834), .b(n1807), .O(n1852));
  andx g1825(.a(n1852), .b(n1331), .O(n1853));
  orx  g1826(.a(n1853), .b(n1851), .O(n1854));
  andx g1827(.a(n1845), .b(n908), .O(n1855));
  andx g1828(.a(n1700), .b(n109), .O(n1856));
  orx  g1829(.a(n1856), .b(n1840), .O(n1857));
  andx g1830(.a(n1857), .b(n228), .O(n1858));
  orx  g1831(.a(n1858), .b(n1855), .O(n1859));
  orx  g1832(.a(n1859), .b(n1854), .O(n1860));
  andx g1833(.a(n1472), .b(n74), .O(n1861));
  andx g1834(.a(n1861), .b(n210), .O(n1862));
  andx g1835(.a(n810), .b(n741), .O(n1863));
  orx  g1836(.a(n1863), .b(n1862), .O(n1864));
  andx g1837(.a(n551), .b(n415), .O(n1865));
  orx  g1838(.a(n1865), .b(n811), .O(n1866));
  orx  g1839(.a(n1866), .b(n1864), .O(n1867));
  andx g1840(.a(n1715), .b(n921), .O(n1868));
  andx g1841(.a(n1827), .b(n974), .O(n1869));
  orx  g1842(.a(n1869), .b(n1868), .O(n1870));
  andx g1843(.a(n1103), .b(n708), .O(n1871));
  andx g1844(.a(n1837), .b(n1331), .O(n1872));
  orx  g1845(.a(n1872), .b(n1871), .O(n1873));
  orx  g1846(.a(n1873), .b(n1870), .O(n1874));
  orx  g1847(.a(n1874), .b(n1867), .O(n1875));
  orx  g1848(.a(n1875), .b(n1860), .O(n1876));
  andx g1849(.a(n1740), .b(n959), .O(n1877));
  andx g1850(.a(n854), .b(n144), .O(n1878));
  andx g1851(.a(n1431), .b(n804), .O(n1879));
  orx  g1852(.a(n1879), .b(n1878), .O(n1880));
  orx  g1853(.a(n1880), .b(n1877), .O(n1881));
  andx g1854(.a(n1749), .b(n551), .O(n1882));
  andx g1855(.a(n1816), .b(n859), .O(n1883));
  orx  g1856(.a(n1883), .b(n1882), .O(n1884));
  orx  g1857(.a(n1884), .b(n1881), .O(n1885));
  andx g1858(.a(n1768), .b(n1056), .O(n1886));
  andx g1859(.a(n1856), .b(n959), .O(n1887));
  orx  g1860(.a(n1887), .b(n1886), .O(n1888));
  orx  g1861(.a(n1431), .b(n759), .O(n1889));
  andx g1862(.a(n1889), .b(n164), .O(n1890));
  orx  g1863(.a(n1890), .b(n761), .O(n1891));
  orx  g1864(.a(n1891), .b(n1888), .O(n1892));
  orx  g1865(.a(n1892), .b(n1885), .O(n1893));
  orx  g1866(.a(n1893), .b(n1876), .O(n1894));
  orx  g1867(.a(n1894), .b(n1850), .O(n1895));
  orx  g1868(.a(n1895), .b(n1802), .O(n1896));
  orx  g1869(.a(n1896), .b(n1785), .O(po05));
  andx g1870(.a(n81), .b(n28), .O(n1898));
  andx g1871(.a(n1898), .b(pi08), .O(n1899));
  andx g1872(.a(n1899), .b(n109), .O(n1900));
  andx g1873(.a(n762), .b(n421), .O(n1901));
  andx g1874(.a(n1471), .b(n421), .O(n1902));
  orx  g1875(.a(n1902), .b(n1901), .O(n1903));
  andx g1876(.a(n1903), .b(n1900), .O(n1904));
  andx g1877(.a(n41), .b(n59), .O(n1905));
  andx g1878(.a(n1905), .b(n36), .O(n1906));
  andx g1879(.a(n1906), .b(n74), .O(n1907));
  andx g1880(.a(n1197), .b(n48), .O(n1908));
  andx g1881(.a(n1908), .b(n910), .O(n1909));
  andx g1882(.a(n1909), .b(n1907), .O(n1910));
  andx g1883(.a(n1910), .b(n28), .O(n1911));
  orx  g1884(.a(n1911), .b(n1904), .O(n1912));
  andx g1885(.a(n60), .b(n276), .O(n1913));
  orx  g1886(.a(n41), .b(pi04), .O(n1914));
  orx  g1887(.a(n1914), .b(n59), .O(n1915));
  invx g1888(.a(n1915), .O(n1916));
  andx g1889(.a(n1916), .b(n1913), .O(n1917));
  andx g1890(.a(n1814), .b(n381), .O(n1918));
  andx g1891(.a(n1918), .b(n31), .O(n1919));
  andx g1892(.a(n1919), .b(n1917), .O(n1920));
  andx g1893(.a(n1917), .b(n1812), .O(n1921));
  andx g1894(.a(n1921), .b(n164), .O(n1922));
  orx  g1895(.a(n1922), .b(n1920), .O(n1923));
  orx  g1896(.a(n1923), .b(n1912), .O(n1924));
  andx g1897(.a(n620), .b(n43), .O(n1925));
  andx g1898(.a(n419), .b(pi07), .O(n1926));
  andx g1899(.a(n1926), .b(n1177), .O(n1927));
  andx g1900(.a(n1927), .b(n1925), .O(n1928));
  andx g1901(.a(n303), .b(n194), .O(n1929));
  andx g1902(.a(n1929), .b(n1902), .O(n1930));
  orx  g1903(.a(n1930), .b(n1928), .O(n1931));
  andx g1904(.a(n327), .b(n77), .O(n1932));
  andx g1905(.a(n1932), .b(n1180), .O(n1933));
  andx g1906(.a(n1933), .b(n1925), .O(n1934));
  andx g1907(.a(n138), .b(n36), .O(n1935));
  andx g1908(.a(n1935), .b(n421), .O(n1936));
  andx g1909(.a(n878), .b(n71), .O(n1937));
  andx g1910(.a(n1937), .b(n209), .O(n1938));
  andx g1911(.a(n1938), .b(n1936), .O(n1939));
  orx  g1912(.a(n1939), .b(n1934), .O(n1940));
  orx  g1913(.a(n1940), .b(n1931), .O(n1941));
  andx g1914(.a(n588), .b(n563), .O(n1942));
  andx g1915(.a(n42), .b(pi04), .O(n1943));
  andx g1916(.a(n1943), .b(n1942), .O(n1944));
  andx g1917(.a(n1944), .b(n1927), .O(n1945));
  andx g1918(.a(n1177), .b(n1015), .O(n1946));
  andx g1919(.a(n1946), .b(n1944), .O(n1947));
  orx  g1920(.a(n1947), .b(n1945), .O(n1948));
  andx g1921(.a(n1937), .b(n361), .O(n1949));
  andx g1922(.a(n1949), .b(n1901), .O(n1950));
  andx g1923(.a(n879), .b(n421), .O(n1951));
  andx g1924(.a(n37), .b(n59), .O(n1952));
  andx g1925(.a(n1952), .b(n36), .O(n1953));
  andx g1926(.a(n1953), .b(n258), .O(n1954));
  andx g1927(.a(n1954), .b(n1951), .O(n1955));
  orx  g1928(.a(n1955), .b(n1950), .O(n1956));
  orx  g1929(.a(n1956), .b(n1948), .O(n1957));
  orx  g1930(.a(n1957), .b(n1941), .O(n1958));
  orx  g1931(.a(n1958), .b(n1924), .O(po06));
  andx g1932(.a(n1944), .b(n1933), .O(n1960));
  orx  g1933(.a(n1960), .b(n1928), .O(n1961));
  andx g1934(.a(n1518), .b(n620), .O(n1962));
  andx g1935(.a(n583), .b(pi07), .O(n1963));
  andx g1936(.a(n1963), .b(n1180), .O(n1964));
  andx g1937(.a(n1964), .b(n1962), .O(n1965));
  orx  g1938(.a(n1965), .b(n1945), .O(n1966));
  orx  g1939(.a(n1966), .b(n1961), .O(n1967));
  andx g1940(.a(n566), .b(n61), .O(n1968));
  andx g1941(.a(n1968), .b(n1814), .O(n1969));
  andx g1942(.a(n1969), .b(n1106), .O(n1970));
  orx  g1943(.a(n1970), .b(n1920), .O(n1971));
  orx  g1944(.a(n1971), .b(n1967), .O(n1972));
  andx g1945(.a(n1953), .b(n71), .O(n1973));
  andx g1946(.a(n910), .b(n74), .O(n1974));
  andx g1947(.a(n1974), .b(n511), .O(n1975));
  andx g1948(.a(n1975), .b(n1973), .O(n1976));
  andx g1949(.a(n1949), .b(n1902), .O(n1977));
  orx  g1950(.a(n1977), .b(n1939), .O(n1978));
  orx  g1951(.a(n1978), .b(n1976), .O(n1979));
  andx g1952(.a(n1935), .b(n258), .O(n1980));
  andx g1953(.a(n240), .b(n90), .O(n1981));
  orx  g1954(.a(n1981), .b(n1980), .O(n1982));
  andx g1955(.a(n1982), .b(n1951), .O(n1983));
  orx  g1956(.a(n1983), .b(n1904), .O(n1984));
  orx  g1957(.a(n1984), .b(n1979), .O(n1985));
  orx  g1958(.a(n1985), .b(n1972), .O(po07));
  orx  g1959(.a(n1594), .b(n1559), .O(n1987));
  andx g1960(.a(n589), .b(n29), .O(n1988));
  andx g1961(.a(n1988), .b(pi12), .O(n1989));
  andx g1962(.a(n1989), .b(n230), .O(n1990));
  andx g1963(.a(n1990), .b(n1987), .O(n1991));
  orx  g1964(.a(n823), .b(n441), .O(n1992));
  andx g1965(.a(n1992), .b(n1989), .O(n1993));
  andx g1966(.a(n680), .b(n109), .O(n1994));
  orx  g1967(.a(n363), .b(n273), .O(n1995));
  orx  g1968(.a(n1995), .b(n1994), .O(n1996));
  andx g1969(.a(n1996), .b(n1056), .O(n1997));
  orx  g1970(.a(n1997), .b(n1993), .O(n1998));
  orx  g1971(.a(n1998), .b(n1991), .O(n1999));
  andx g1972(.a(n1913), .b(n224), .O(n2000));
  andx g1973(.a(n961), .b(n224), .O(n2001));
  orx  g1974(.a(n2001), .b(n2000), .O(n2002));
  andx g1975(.a(n1812), .b(n1271), .O(n2003));
  andx g1976(.a(n2003), .b(n1907), .O(n2004));
  orx  g1977(.a(n2004), .b(n1208), .O(n2005));
  orx  g1978(.a(n2005), .b(n2002), .O(n2006));
  andx g1979(.a(n565), .b(n265), .O(n2007));
  andx g1980(.a(n1899), .b(n240), .O(n2008));
  andx g1981(.a(n2008), .b(n1936), .O(n2009));
  orx  g1982(.a(n2009), .b(n2007), .O(n2010));
  andx g1983(.a(n565), .b(n267), .O(n2011));
  andx g1984(.a(n957), .b(n292), .O(n2012));
  orx  g1985(.a(n2012), .b(n2011), .O(n2013));
  orx  g1986(.a(n2013), .b(n2010), .O(n2014));
  orx  g1987(.a(n2014), .b(n2006), .O(n2015));
  andx g1988(.a(n1065), .b(n688), .O(n2016));
  andx g1989(.a(n1065), .b(n669), .O(n2017));
  andx g1990(.a(n1056), .b(n155), .O(n2018));
  andx g1991(.a(n133), .b(pi03), .O(n2019));
  andx g1992(.a(n2019), .b(n61), .O(n2020));
  andx g1993(.a(n2020), .b(n132), .O(n2021));
  orx  g1994(.a(n2021), .b(n2018), .O(n2022));
  orx  g1995(.a(n2022), .b(n2017), .O(n2023));
  orx  g1996(.a(n2023), .b(n2016), .O(n2024));
  orx  g1997(.a(n2024), .b(n2015), .O(n2025));
  orx  g1998(.a(n2025), .b(n1999), .O(n2026));
  andx g1999(.a(n1913), .b(n29), .O(n2027));
  orx  g2000(.a(n1667), .b(n669), .O(n2028));
  orx  g2001(.a(n2028), .b(n689), .O(n2029));
  andx g2002(.a(n2029), .b(n2027), .O(n2030));
  andx g2003(.a(n1592), .b(n30), .O(n2031));
  orx  g2004(.a(n203), .b(n164), .O(n2032));
  orx  g2005(.a(n340), .b(n124), .O(n2033));
  orx  g2006(.a(n2033), .b(n2032), .O(n2034));
  orx  g2007(.a(n2034), .b(n2031), .O(n2035));
  andx g2008(.a(n61), .b(pi03), .O(n2036));
  andx g2009(.a(n2036), .b(n42), .O(n2037));
  andx g2010(.a(n2037), .b(n2035), .O(n2038));
  orx  g2011(.a(n2038), .b(n2030), .O(n2039));
  orx  g2012(.a(n2039), .b(n2026), .O(n2040));
  andx g2013(.a(n1512), .b(n822), .O(n2041));
  orx  g2014(.a(n2041), .b(n1574), .O(n2042));
  orx  g2015(.a(n2042), .b(n1578), .O(n2043));
  andx g2016(.a(n2043), .b(pi12), .O(n2044));
  orx  g2017(.a(n671), .b(n637), .O(n2045));
  andx g2018(.a(n1512), .b(pi12), .O(n2046));
  andx g2019(.a(n2046), .b(n1594), .O(n2047));
  orx  g2020(.a(n2047), .b(n667), .O(n2048));
  orx  g2021(.a(n2048), .b(n2045), .O(n2049));
  orx  g2022(.a(n2049), .b(n2044), .O(n2050));
  andx g2023(.a(n2050), .b(n2027), .O(n2051));
  andx g2024(.a(n1622), .b(n741), .O(n2052));
  orx  g2025(.a(n2052), .b(n1886), .O(n2053));
  andx g2026(.a(n2045), .b(n1065), .O(n2054));
  andx g2027(.a(n1620), .b(n741), .O(n2055));
  orx  g2028(.a(n2055), .b(n2054), .O(n2056));
  orx  g2029(.a(n2056), .b(n2053), .O(n2057));
  andx g2030(.a(n1056), .b(n149), .O(n2058));
  orx  g2031(.a(n2058), .b(n1910), .O(n2059));
  orx  g2032(.a(n1879), .b(n1681), .O(n2060));
  orx  g2033(.a(n2060), .b(n2059), .O(n2061));
  andx g2034(.a(n2036), .b(n292), .O(n2062));
  andx g2035(.a(n2020), .b(n69), .O(n2063));
  orx  g2036(.a(n2063), .b(n2062), .O(n2064));
  andx g2037(.a(n1913), .b(n695), .O(n2065));
  orx  g2038(.a(n2065), .b(n1939), .O(n2066));
  orx  g2039(.a(n2066), .b(n2064), .O(n2067));
  orx  g2040(.a(n2067), .b(n2061), .O(n2068));
  orx  g2041(.a(n2068), .b(n2057), .O(n2069));
  andx g2042(.a(n1618), .b(n741), .O(n2070));
  andx g2043(.a(n1988), .b(n738), .O(n2071));
  orx  g2044(.a(n2071), .b(n1092), .O(n2072));
  andx g2045(.a(n1084), .b(n741), .O(n2073));
  andx g2046(.a(n957), .b(n484), .O(n2074));
  orx  g2047(.a(n2074), .b(n1757), .O(n2075));
  orx  g2048(.a(n2075), .b(n2073), .O(n2076));
  orx  g2049(.a(n2076), .b(n2072), .O(n2077));
  orx  g2050(.a(n2077), .b(n2070), .O(n2078));
  orx  g2051(.a(n2078), .b(n2069), .O(n2079));
  orx  g2052(.a(n2079), .b(n2051), .O(n2080));
  orx  g2053(.a(n2080), .b(n2040), .O(po08));
  andx g2054(.a(n1565), .b(n896), .O(n2082));
  andx g2055(.a(n1943), .b(n1593), .O(n2083));
  orx  g2056(.a(n2083), .b(n2016), .O(n2084));
  orx  g2057(.a(n1577), .b(n128), .O(n2085));
  orx  g2058(.a(n2085), .b(n2084), .O(n2086));
  andx g2059(.a(n1942), .b(n316), .O(n2087));
  andx g2060(.a(n853), .b(n484), .O(n2088));
  andx g2061(.a(n89), .b(pi01), .O(n2089));
  andx g2062(.a(n2089), .b(pi13), .O(n2090));
  andx g2063(.a(n2090), .b(n112), .O(n2091));
  orx  g2064(.a(n2091), .b(n2088), .O(n2092));
  orx  g2065(.a(n2092), .b(n2087), .O(n2093));
  orx  g2066(.a(n2093), .b(n55), .O(n2094));
  andx g2067(.a(n1996), .b(n854), .O(n2095));
  andx g2068(.a(n81), .b(n77), .O(n2096));
  andx g2069(.a(n2096), .b(n101), .O(n2097));
  andx g2070(.a(n2097), .b(n327), .O(n2098));
  andx g2071(.a(n2098), .b(n1962), .O(n2099));
  orx  g2072(.a(n2099), .b(n1934), .O(n2100));
  orx  g2073(.a(n2100), .b(n2095), .O(n2101));
  orx  g2074(.a(n2101), .b(n2094), .O(n2102));
  orx  g2075(.a(n2102), .b(n2086), .O(n2103));
  orx  g2076(.a(n2103), .b(n2082), .O(n2104));
  andx g2077(.a(n1547), .b(n896), .O(n2105));
  andx g2078(.a(n1942), .b(n100), .O(n2106));
  andx g2079(.a(n2106), .b(n390), .O(n2107));
  orx  g2080(.a(n2107), .b(n2105), .O(n2108));
  andx g2081(.a(n1611), .b(n254), .O(n2109));
  andx g2082(.a(n1035), .b(n312), .O(n2110));
  orx  g2083(.a(n2110), .b(n2109), .O(n2111));
  orx  g2084(.a(n2111), .b(n2108), .O(n2112));
  andx g2085(.a(n1943), .b(n565), .O(n2113));
  andx g2086(.a(n2113), .b(n203), .O(n2114));
  andx g2087(.a(n1035), .b(n413), .O(n2115));
  orx  g2088(.a(n2115), .b(n2114), .O(n2116));
  andx g2089(.a(n1901), .b(n1900), .O(n2117));
  andx g2090(.a(n1547), .b(n576), .O(n2118));
  orx  g2091(.a(n2118), .b(n2117), .O(n2119));
  orx  g2092(.a(n2119), .b(n2116), .O(n2120));
  orx  g2093(.a(n2120), .b(n2112), .O(n2121));
  andx g2094(.a(n1036), .b(n547), .O(n2122));
  orx  g2095(.a(n2122), .b(n1202), .O(n2123));
  andx g2096(.a(n385), .b(pi02), .O(n2124));
  andx g2097(.a(n2124), .b(n182), .O(n2125));
  andx g2098(.a(n2125), .b(n2090), .O(n2126));
  orx  g2099(.a(n2126), .b(n552), .O(n2127));
  orx  g2100(.a(n2127), .b(n2123), .O(n2128));
  andx g2101(.a(n2113), .b(n340), .O(n2129));
  andx g2102(.a(n1518), .b(n565), .O(n2130));
  andx g2103(.a(n2130), .b(n203), .O(n2131));
  orx  g2104(.a(n2131), .b(n2129), .O(n2132));
  andx g2105(.a(n133), .b(pi04), .O(n2133));
  andx g2106(.a(n2133), .b(n565), .O(n2134));
  andx g2107(.a(n2134), .b(n132), .O(n2135));
  andx g2108(.a(n2130), .b(n340), .O(n2136));
  orx  g2109(.a(n2136), .b(n2135), .O(n2137));
  orx  g2110(.a(n2137), .b(n2132), .O(n2138));
  orx  g2111(.a(n2138), .b(n2128), .O(n2139));
  orx  g2112(.a(n2139), .b(n2121), .O(n2140));
  orx  g2113(.a(n1724), .b(n1681), .O(n2141));
  andx g2114(.a(n854), .b(n149), .O(n2142));
  orx  g2115(.a(n2142), .b(n1216), .O(n2143));
  orx  g2116(.a(n2143), .b(n2141), .O(n2144));
  andx g2117(.a(n1518), .b(n837), .O(n2145));
  orx  g2118(.a(n2145), .b(n1557), .O(n2146));
  andx g2119(.a(n2146), .b(n576), .O(n2147));
  andx g2120(.a(n2113), .b(n124), .O(n2148));
  orx  g2121(.a(n2148), .b(n2147), .O(n2149));
  orx  g2122(.a(n2149), .b(n2144), .O(n2150));
  orx  g2123(.a(n1977), .b(n1757), .O(n2151));
  andx g2124(.a(n2090), .b(n115), .O(n2152));
  orx  g2125(.a(n2152), .b(n1955), .O(n2153));
  orx  g2126(.a(n2153), .b(n2151), .O(n2154));
  andx g2127(.a(n172), .b(n2130), .O(n2155));
  orx  g2128(.a(n2155), .b(n2001), .O(n2156));
  andx g2129(.a(n853), .b(n292), .O(n2157));
  andx g2130(.a(n2113), .b(n164), .O(n2158));
  orx  g2131(.a(n2158), .b(n2157), .O(n2159));
  orx  g2132(.a(n2159), .b(n2156), .O(n2160));
  orx  g2133(.a(n2160), .b(n2154), .O(n2161));
  orx  g2134(.a(n2161), .b(n2150), .O(n2162));
  orx  g2135(.a(n2162), .b(n2140), .O(n2163));
  andx g2136(.a(n1035), .b(n348), .O(n2164));
  andx g2137(.a(n180), .b(n32), .O(n2165));
  andx g2138(.a(n2165), .b(n393), .O(n2166));
  orx  g2139(.a(n2166), .b(n2164), .O(n2167));
  orx  g2140(.a(n352), .b(n317), .O(n2168));
  orx  g2141(.a(n2168), .b(n2167), .O(n2169));
  andx g2142(.a(n685), .b(pi13), .O(n2170));
  andx g2143(.a(n2170), .b(n828), .O(n2171));
  andx g2144(.a(n1035), .b(n402), .O(n2172));
  orx  g2145(.a(n2172), .b(n2171), .O(n2173));
  orx  g2146(.a(n1112), .b(n507), .O(n2174));
  orx  g2147(.a(n2174), .b(n2173), .O(n2175));
  orx  g2148(.a(n2175), .b(n2169), .O(n2176));
  andx g2149(.a(n1524), .b(n896), .O(n2177));
  orx  g2150(.a(n2177), .b(n384), .O(n2178));
  andx g2151(.a(n685), .b(n620), .O(n2179));
  andx g2152(.a(n2179), .b(n515), .O(n2180));
  orx  g2153(.a(n2180), .b(n238), .O(n2181));
  orx  g2154(.a(n2181), .b(n2178), .O(n2182));
  andx g2155(.a(n69), .b(n58), .O(n2183));
  orx  g2156(.a(n2183), .b(n429), .O(n2184));
  orx  g2157(.a(n2017), .b(n1550), .O(n2185));
  orx  g2158(.a(n2185), .b(n2184), .O(n2186));
  orx  g2159(.a(n2186), .b(n2182), .O(n2187));
  orx  g2160(.a(n2187), .b(n2176), .O(n2188));
  orx  g2161(.a(n539), .b(n418), .O(n2189));
  orx  g2162(.a(n1090), .b(n855), .O(n2190));
  orx  g2163(.a(n2190), .b(n2189), .O(n2191));
  andx g2164(.a(n1942), .b(n103), .O(n2192));
  andx g2165(.a(n2192), .b(n1568), .O(n2193));
  orx  g2166(.a(n2193), .b(n1514), .O(n2194));
  orx  g2167(.a(n2009), .b(n1976), .O(n2195));
  orx  g2168(.a(n2195), .b(n2194), .O(n2196));
  orx  g2169(.a(n2196), .b(n2191), .O(n2197));
  andx g2170(.a(n854), .b(n155), .O(n2198));
  orx  g2171(.a(n2198), .b(n377), .O(n2199));
  andx g2172(.a(n2090), .b(n520), .O(n2200));
  orx  g2173(.a(n2200), .b(n936), .O(n2201));
  orx  g2174(.a(n2201), .b(n2199), .O(n2202));
  andx g2175(.a(n2179), .b(n104), .O(n2203));
  orx  g2176(.a(n2203), .b(n449), .O(n2204));
  andx g2177(.a(n2170), .b(n827), .O(n2205));
  orx  g2178(.a(n2205), .b(n606), .O(n2206));
  orx  g2179(.a(n2206), .b(n2204), .O(n2207));
  orx  g2180(.a(n2207), .b(n2202), .O(n2208));
  orx  g2181(.a(n2208), .b(n2197), .O(n2209));
  orx  g2182(.a(n2209), .b(n2188), .O(n2210));
  orx  g2183(.a(n2210), .b(n2163), .O(n2211));
  andx g2184(.a(n1942), .b(pi13), .O(n2212));
  orx  g2185(.a(n1761), .b(n359), .O(n2213));
  andx g2186(.a(n2213), .b(n2212), .O(n2214));
  orx  g2187(.a(n494), .b(n372), .O(n2215));
  andx g2188(.a(n2215), .b(n2090), .O(n2216));
  andx g2189(.a(n1584), .b(n254), .O(n2217));
  andx g2190(.a(n1512), .b(n1500), .O(n2218));
  andx g2191(.a(n2218), .b(n1062), .O(n2219));
  orx  g2192(.a(n2219), .b(n2217), .O(n2220));
  orx  g2193(.a(n2220), .b(n2216), .O(n2221));
  orx  g2194(.a(n2221), .b(n2214), .O(n2222));
  orx  g2195(.a(n2222), .b(n544), .O(n2223));
  orx  g2196(.a(n2054), .b(n1880), .O(n2224));
  orx  g2197(.a(n550), .b(n183), .O(n2225));
  andx g2198(.a(n2225), .b(n2212), .O(n2226));
  andx g2199(.a(n209), .b(n90), .O(n2227));
  andx g2200(.a(n297), .b(n122), .O(n2228));
  andx g2201(.a(n2228), .b(n2227), .O(n2229));
  orx  g2202(.a(n2229), .b(n1950), .O(n2230));
  orx  g2203(.a(n2230), .b(n2226), .O(n2231));
  orx  g2204(.a(n2231), .b(n2224), .O(n2232));
  orx  g2205(.a(n1567), .b(n428), .O(n2233));
  andx g2206(.a(n2233), .b(n1942), .O(n2234));
  andx g2207(.a(n1790), .b(n254), .O(n2235));
  orx  g2208(.a(n2235), .b(n400), .O(n2236));
  orx  g2209(.a(n2236), .b(n2234), .O(n2237));
  andx g2210(.a(n1558), .b(n1512), .O(n2238));
  andx g2211(.a(n2238), .b(n1062), .O(n2239));
  orx  g2212(.a(n2239), .b(n342), .O(n2240));
  orx  g2213(.a(n2240), .b(n2237), .O(n2241));
  orx  g2214(.a(n2241), .b(n2232), .O(n2242));
  andx g2215(.a(n1518), .b(n750), .O(n2243));
  andx g2216(.a(n2243), .b(n576), .O(n2244));
  andx g2217(.a(n2032), .b(n45), .O(n2245));
  orx  g2218(.a(n2245), .b(n2244), .O(n2246));
  orx  g2219(.a(n2124), .b(n361), .O(n2247));
  andx g2220(.a(n2247), .b(n2089), .O(n2248));
  andx g2221(.a(n2248), .b(n217), .O(n2249));
  orx  g2222(.a(n2249), .b(n1668), .O(n2250));
  orx  g2223(.a(n2250), .b(n2246), .O(n2251));
  orx  g2224(.a(n1961), .b(n768), .O(n2252));
  andx g2225(.a(n1655), .b(n701), .O(n2253));
  andx g2226(.a(n696), .b(n565), .O(n2254));
  orx  g2227(.a(n2254), .b(n2253), .O(n2255));
  orx  g2228(.a(n2255), .b(n2252), .O(n2256));
  orx  g2229(.a(n2256), .b(n2251), .O(n2257));
  orx  g2230(.a(n2257), .b(n2242), .O(n2258));
  orx  g2231(.a(n2258), .b(n2223), .O(n2259));
  orx  g2232(.a(n2259), .b(n2211), .O(n2260));
  orx  g2233(.a(n2260), .b(n2104), .O(po09));
  andx g2234(.a(n122), .b(n109), .O(n2262));
  orx  g2235(.a(n2262), .b(n1281), .O(n2263));
  andx g2236(.a(n1179), .b(pi08), .O(n2264));
  andx g2237(.a(n2264), .b(n361), .O(n2265));
  andx g2238(.a(n1271), .b(n152), .O(n2266));
  orx  g2239(.a(n2266), .b(n2265), .O(n2267));
  orx  g2240(.a(n2267), .b(n2263), .O(n2268));
  andx g2241(.a(n2268), .b(n228), .O(n2269));
  andx g2242(.a(n896), .b(n704), .O(n2270));
  andx g2243(.a(n921), .b(n786), .O(n2271));
  orx  g2244(.a(n2271), .b(n2270), .O(n2272));
  andx g2245(.a(n2272), .b(n1271), .O(n2273));
  orx  g2246(.a(n2273), .b(n2269), .O(n2274));
  andx g2247(.a(n240), .b(n122), .O(n2275));
  andx g2248(.a(n2275), .b(n1347), .O(n2276));
  andx g2249(.a(n2262), .b(n958), .O(n2277));
  orx  g2250(.a(n2277), .b(n898), .O(n2278));
  orx  g2251(.a(n2278), .b(n2276), .O(n2279));
  orx  g2252(.a(n2279), .b(n966), .O(n2280));
  orx  g2253(.a(n2280), .b(n2274), .O(n2281));
  andx g2254(.a(n942), .b(n480), .O(n2282));
  andx g2255(.a(n2282), .b(n278), .O(n2283));
  orx  g2256(.a(n2283), .b(n1490), .O(n2284));
  andx g2257(.a(n406), .b(n146), .O(n2285));
  andx g2258(.a(n2285), .b(n278), .O(n2286));
  orx  g2259(.a(n2286), .b(n169), .O(n2287));
  orx  g2260(.a(n2287), .b(n2284), .O(n2288));
  andx g2261(.a(n1790), .b(n178), .O(n2289));
  andx g2262(.a(n2265), .b(n956), .O(n2290));
  orx  g2263(.a(n2290), .b(n2289), .O(n2291));
  orx  g2264(.a(n2172), .b(n403), .O(n2292));
  orx  g2265(.a(n2292), .b(n2291), .O(n2293));
  orx  g2266(.a(n2293), .b(n2288), .O(n2294));
  orx  g2267(.a(n2282), .b(n857), .O(n2295));
  andx g2268(.a(n2295), .b(n859), .O(n2296));
  orx  g2269(.a(n2296), .b(n1064), .O(n2297));
  andx g2270(.a(n1065), .b(n671), .O(n2298));
  andx g2271(.a(n908), .b(n789), .O(n2299));
  orx  g2272(.a(n2299), .b(n2298), .O(n2300));
  andx g2273(.a(n908), .b(n756), .O(n2301));
  orx  g2274(.a(n2301), .b(n2058), .O(n2302));
  orx  g2275(.a(n2302), .b(n2300), .O(n2303));
  orx  g2276(.a(n2303), .b(n2297), .O(n2304));
  orx  g2277(.a(n2304), .b(n2294), .O(n2305));
  orx  g2278(.a(n2305), .b(n2281), .O(n2306));
  andx g2279(.a(n1814), .b(n242), .O(n2307));
  orx  g2280(.a(n1097), .b(n239), .O(n2308));
  orx  g2281(.a(n2308), .b(n1040), .O(n2309));
  andx g2282(.a(n2309), .b(n2307), .O(n2310));
  orx  g2283(.a(n1356), .b(n548), .O(n2311));
  andx g2284(.a(n1812), .b(n242), .O(n2312));
  andx g2285(.a(n2312), .b(n2311), .O(n2313));
  orx  g2286(.a(n1035), .b(n858), .O(n2314));
  andx g2287(.a(n1811), .b(n166), .O(n2315));
  andx g2288(.a(n2315), .b(n2314), .O(n2316));
  andx g2289(.a(n2316), .b(n492), .O(n2317));
  andx g2290(.a(n1963), .b(n872), .O(n2318));
  andx g2291(.a(n2318), .b(n1243), .O(n2319));
  orx  g2292(.a(n2319), .b(n2317), .O(n2320));
  orx  g2293(.a(n2320), .b(n2313), .O(n2321));
  orx  g2294(.a(n2321), .b(n2310), .O(n2322));
  andx g2295(.a(n2264), .b(n209), .O(n2323));
  orx  g2296(.a(n2323), .b(n1264), .O(n2324));
  andx g2297(.a(n1271), .b(n786), .O(n2325));
  orx  g2298(.a(n2325), .b(n2275), .O(n2326));
  orx  g2299(.a(n2326), .b(n2324), .O(n2327));
  andx g2300(.a(n2327), .b(n1062), .O(n2328));
  orx  g2301(.a(n2328), .b(n973), .O(n2329));
  andx g2302(.a(n231), .b(n209), .O(n2330));
  orx  g2303(.a(n2330), .b(n912), .O(n2331));
  orx  g2304(.a(n2331), .b(n2324), .O(n2332));
  andx g2305(.a(n2332), .b(n909), .O(n2333));
  orx  g2306(.a(n2330), .b(n850), .O(n2334));
  orx  g2307(.a(n2334), .b(n2324), .O(n2335));
  andx g2308(.a(n2335), .b(n576), .O(n2336));
  orx  g2309(.a(n2336), .b(n2333), .O(n2337));
  orx  g2310(.a(n2337), .b(n2329), .O(n2338));
  orx  g2311(.a(n2338), .b(n2322), .O(n2339));
  orx  g2312(.a(n2339), .b(n2306), .O(n2340));
  andx g2313(.a(n1281), .b(n959), .O(n2341));
  andx g2314(.a(n1194), .b(n328), .O(n2342));
  andx g2315(.a(n1194), .b(n406), .O(n2343));
  orx  g2316(.a(n2343), .b(n2342), .O(n2344));
  andx g2317(.a(n2344), .b(n859), .O(n2345));
  orx  g2318(.a(n2345), .b(n2341), .O(n2346));
  orx  g2319(.a(n789), .b(n756), .O(n2347));
  andx g2320(.a(n2347), .b(n1103), .O(n2348));
  orx  g2321(.a(n2348), .b(n1052), .O(n2349));
  orx  g2322(.a(n2349), .b(n2346), .O(n2350));
  andx g2323(.a(n2347), .b(n741), .O(n2351));
  orx  g2324(.a(n2342), .b(n857), .O(n2352));
  andx g2325(.a(n2352), .b(n278), .O(n2353));
  orx  g2326(.a(n2353), .b(n2351), .O(n2354));
  andx g2327(.a(n150), .b(n47), .O(n2355));
  andx g2328(.a(n2262), .b(n956), .O(n2356));
  andx g2329(.a(n962), .b(n123), .O(n2357));
  orx  g2330(.a(n2357), .b(n2356), .O(n2358));
  orx  g2331(.a(n2358), .b(n2355), .O(n2359));
  orx  g2332(.a(n2359), .b(n2354), .O(n2360));
  orx  g2333(.a(n2360), .b(n2350), .O(n2361));
  andx g2334(.a(n1387), .b(n86), .O(n2362));
  orx  g2335(.a(n2362), .b(n914), .O(n2363));
  andx g2336(.a(n2363), .b(n586), .O(n2364));
  andx g2337(.a(n2318), .b(n1010), .O(n2365));
  andx g2338(.a(n1963), .b(n502), .O(n2366));
  andx g2339(.a(n2366), .b(n914), .O(n2367));
  orx  g2340(.a(n2367), .b(n2365), .O(n2368));
  andx g2341(.a(n2324), .b(n921), .O(n2369));
  orx  g2342(.a(n2369), .b(n2368), .O(n2370));
  andx g2343(.a(n30), .b(pi08), .O(n2371));
  andx g2344(.a(n2371), .b(n1179), .O(n2372));
  andx g2345(.a(n2372), .b(n996), .O(n2373));
  andx g2346(.a(n2347), .b(n1020), .O(n2374));
  orx  g2347(.a(n2374), .b(n2373), .O(n2375));
  orx  g2348(.a(n2375), .b(n2370), .O(n2376));
  orx  g2349(.a(n2376), .b(n2364), .O(n2377));
  orx  g2350(.a(n2377), .b(n2361), .O(n2378));
  andx g2351(.a(n1390), .b(n344), .O(n2379));
  orx  g2352(.a(n2379), .b(n1880), .O(n2380));
  andx g2353(.a(n2372), .b(n993), .O(n2381));
  orx  g2354(.a(n2343), .b(n1293), .O(n2382));
  andx g2355(.a(n2382), .b(n278), .O(n2383));
  orx  g2356(.a(n2383), .b(n2381), .O(n2384));
  orx  g2357(.a(n2384), .b(n2380), .O(n2385));
  andx g2358(.a(n2307), .b(n941), .O(n2386));
  orx  g2359(.a(n2386), .b(n866), .O(n2387));
  orx  g2360(.a(n2330), .b(n2325), .O(n2388));
  andx g2361(.a(n2388), .b(n896), .O(n2389));
  orx  g2362(.a(n2389), .b(n2387), .O(n2390));
  andx g2363(.a(n2326), .b(n909), .O(n2391));
  andx g2364(.a(n2347), .b(n701), .O(n2392));
  orx  g2365(.a(n2392), .b(n2391), .O(n2393));
  orx  g2366(.a(n2393), .b(n2390), .O(n2394));
  orx  g2367(.a(n2394), .b(n2385), .O(n2395));
  andx g2368(.a(n1796), .b(n858), .O(n2396));
  andx g2369(.a(n1852), .b(n871), .O(n2397));
  orx  g2370(.a(n2397), .b(n2396), .O(n2398));
  andx g2371(.a(n2326), .b(n576), .O(n2399));
  orx  g2372(.a(n2399), .b(n353), .O(n2400));
  orx  g2373(.a(n2400), .b(n2398), .O(n2401));
  andx g2374(.a(n2266), .b(n959), .O(n2402));
  orx  g2375(.a(n2402), .b(n2236), .O(n2403));
  orx  g2376(.a(n1142), .b(n979), .O(n2404));
  orx  g2377(.a(n2404), .b(n2403), .O(n2405));
  orx  g2378(.a(n2405), .b(n2401), .O(n2406));
  orx  g2379(.a(n2406), .b(n2395), .O(n2407));
  andx g2380(.a(n172), .b(n574), .O(n2408));
  andx g2381(.a(n1056), .b(n144), .O(n2409));
  orx  g2382(.a(n2409), .b(n2408), .O(n2410));
  orx  g2383(.a(n2142), .b(n805), .O(n2411));
  orx  g2384(.a(n2411), .b(n2410), .O(n2412));
  andx g2385(.a(n1611), .b(n139), .O(n2413));
  andx g2386(.a(n1271), .b(n668), .O(n2414));
  andx g2387(.a(n2414), .b(n1523), .O(n2415));
  orx  g2388(.a(n2415), .b(n2413), .O(n2416));
  andx g2389(.a(n2330), .b(n1062), .O(n2417));
  andx g2390(.a(n361), .b(n231), .O(n2418));
  andx g2391(.a(n2418), .b(n228), .O(n2419));
  orx  g2392(.a(n2419), .b(n2417), .O(n2420));
  orx  g2393(.a(n2420), .b(n2416), .O(n2421));
  orx  g2394(.a(n2421), .b(n2412), .O(n2422));
  andx g2395(.a(n1355), .b(n348), .O(n2423));
  andx g2396(.a(n2418), .b(n956), .O(n2424));
  orx  g2397(.a(n2424), .b(n2423), .O(n2425));
  andx g2398(.a(n974), .b(n123), .O(n2426));
  orx  g2399(.a(n2426), .b(n975), .O(n2427));
  orx  g2400(.a(n2427), .b(n2425), .O(n2428));
  orx  g2401(.a(n1443), .b(n1235), .O(n2429));
  andx g2402(.a(n2330), .b(n921), .O(n2430));
  orx  g2403(.a(n2430), .b(n587), .O(n2431));
  orx  g2404(.a(n2431), .b(n2429), .O(n2432));
  orx  g2405(.a(n2432), .b(n2428), .O(n2433));
  orx  g2406(.a(n2433), .b(n2422), .O(n2434));
  andx g2407(.a(n1790), .b(n940), .O(n2435));
  orx  g2408(.a(n2435), .b(n1495), .O(n2436));
  andx g2409(.a(n858), .b(n334), .O(n2437));
  andx g2410(.a(n2307), .b(n1078), .O(n2438));
  orx  g2411(.a(n2438), .b(n2437), .O(n2439));
  orx  g2412(.a(n2439), .b(n2436), .O(n2440));
  orx  g2413(.a(n2285), .b(n1293), .O(n2441));
  andx g2414(.a(n2441), .b(n859), .O(n2442));
  andx g2415(.a(n608), .b(n76), .O(n2443));
  orx  g2416(.a(n2443), .b(n2109), .O(n2444));
  orx  g2417(.a(n2444), .b(n2442), .O(n2445));
  orx  g2418(.a(n2445), .b(n2440), .O(n2446));
  andx g2419(.a(n1331), .b(n76), .O(n2447));
  andx g2420(.a(n473), .b(n323), .O(n2448));
  orx  g2421(.a(n2448), .b(n2447), .O(n2449));
  andx g2422(.a(n995), .b(n344), .O(n2450));
  andx g2423(.a(n1611), .b(n940), .O(n2451));
  orx  g2424(.a(n2451), .b(n2450), .O(n2452));
  orx  g2425(.a(n2452), .b(n2449), .O(n2453));
  orx  g2426(.a(n858), .b(n178), .O(n2454));
  andx g2427(.a(n2454), .b(n1611), .O(n2455));
  orx  g2428(.a(n2455), .b(n366), .O(n2456));
  andx g2429(.a(n2366), .b(n581), .O(n2457));
  andx g2430(.a(n402), .b(n95), .O(n2458));
  orx  g2431(.a(n2458), .b(n2457), .O(n2459));
  orx  g2432(.a(n2459), .b(n2456), .O(n2460));
  orx  g2433(.a(n2460), .b(n2453), .O(n2461));
  orx  g2434(.a(n2461), .b(n2446), .O(n2462));
  orx  g2435(.a(n2462), .b(n2434), .O(n2463));
  orx  g2436(.a(n2463), .b(n2407), .O(n2464));
  orx  g2437(.a(n2464), .b(n2378), .O(n2465));
  orx  g2438(.a(n2465), .b(n2340), .O(po10));
  orx  g2439(.a(n1054), .b(n57), .O(n2467));
  andx g2440(.a(n2467), .b(n267), .O(n2468));
  andx g2441(.a(n533), .b(n71), .O(n2469));
  andx g2442(.a(n2469), .b(n193), .O(n2470));
  andx g2443(.a(n109), .b(n35), .O(n2471));
  orx  g2444(.a(n2471), .b(n974), .O(n2472));
  orx  g2445(.a(n2472), .b(n964), .O(n2473));
  andx g2446(.a(n2473), .b(n2470), .O(n2474));
  orx  g2447(.a(n2474), .b(n2468), .O(n2475));
  orx  g2448(.a(n2297), .b(n2279), .O(n2476));
  orx  g2449(.a(n2476), .b(n2475), .O(n2477));
  orx  g2450(.a(n2477), .b(n2322), .O(n2478));
  orx  g2451(.a(n2478), .b(n982), .O(n2479));
  orx  g2452(.a(n974), .b(n962), .O(n2480));
  andx g2453(.a(n2480), .b(n33), .O(n2481));
  orx  g2454(.a(n2481), .b(n326), .O(n2482));
  andx g2455(.a(n2470), .b(n109), .O(n2483));
  andx g2456(.a(n2483), .b(n959), .O(n2484));
  andx g2457(.a(n534), .b(n240), .O(n2485));
  orx  g2458(.a(n2485), .b(n2275), .O(n2486));
  andx g2459(.a(n2486), .b(n909), .O(n2487));
  orx  g2460(.a(n2487), .b(n2484), .O(n2488));
  orx  g2461(.a(n2488), .b(n2482), .O(n2489));
  andx g2462(.a(n2470), .b(n240), .O(n2490));
  andx g2463(.a(n2490), .b(n1537), .O(n2491));
  orx  g2464(.a(n2491), .b(n1142), .O(n2492));
  orx  g2465(.a(n2075), .b(n318), .O(n2493));
  orx  g2466(.a(n2493), .b(n2492), .O(n2494));
  orx  g2467(.a(n2494), .b(n2489), .O(n2495));
  andx g2468(.a(n1814), .b(n283), .O(n2496));
  orx  g2469(.a(n2308), .b(n1078), .O(n2497));
  andx g2470(.a(n2497), .b(n2496), .O(n2498));
  andx g2471(.a(n2490), .b(n1073), .O(n2499));
  andx g2472(.a(n1494), .b(n146), .O(n2500));
  andx g2473(.a(n2500), .b(n1057), .O(n2501));
  orx  g2474(.a(n2501), .b(n2499), .O(n2502));
  orx  g2475(.a(n1040), .b(n941), .O(n2503));
  andx g2476(.a(n2503), .b(n2496), .O(n2504));
  orx  g2477(.a(n2504), .b(n2387), .O(n2505));
  orx  g2478(.a(n2505), .b(n2502), .O(n2506));
  orx  g2479(.a(n2506), .b(n2498), .O(n2507));
  orx  g2480(.a(n2507), .b(n2495), .O(n2508));
  andx g2481(.a(n484), .b(n35), .O(n2509));
  andx g2482(.a(n657), .b(n119), .O(n2510));
  andx g2483(.a(n2510), .b(n323), .O(n2511));
  orx  g2484(.a(n2511), .b(n2509), .O(n2512));
  orx  g2485(.a(n2438), .b(n1477), .O(n2513));
  orx  g2486(.a(n2513), .b(n2512), .O(n2514));
  andx g2487(.a(n1812), .b(n283), .O(n2515));
  andx g2488(.a(n2515), .b(n1037), .O(n2516));
  orx  g2489(.a(n2516), .b(n2368), .O(n2517));
  orx  g2490(.a(n2517), .b(n2514), .O(n2518));
  andx g2491(.a(n1328), .b(n942), .O(n2519));
  andx g2492(.a(n323), .b(n30), .O(n2520));
  andx g2493(.a(n2520), .b(n2519), .O(n2521));
  andx g2494(.a(n1010), .b(n79), .O(n2522));
  orx  g2495(.a(n2522), .b(n2521), .O(n2523));
  orx  g2496(.a(n2523), .b(n1052), .O(n2524));
  andx g2497(.a(n1070), .b(n79), .O(n2525));
  andx g2498(.a(n963), .b(n33), .O(n2526));
  orx  g2499(.a(n2526), .b(n2525), .O(n2527));
  andx g2500(.a(n858), .b(n69), .O(n2528));
  orx  g2501(.a(n2528), .b(n809), .O(n2529));
  orx  g2502(.a(n2529), .b(n2527), .O(n2530));
  orx  g2503(.a(n2530), .b(n2524), .O(n2531));
  orx  g2504(.a(n2531), .b(n2518), .O(n2532));
  andx g2505(.a(n2316), .b(n515), .O(n2533));
  orx  g2506(.a(n2533), .b(n2358), .O(n2534));
  andx g2507(.a(n398), .b(n146), .O(n2535));
  andx g2508(.a(n2535), .b(n1026), .O(n2536));
  andx g2509(.a(n2535), .b(n1338), .O(n2537));
  orx  g2510(.a(n2537), .b(n2536), .O(n2538));
  orx  g2511(.a(n2538), .b(n2534), .O(n2539));
  andx g2512(.a(n1814), .b(n143), .O(n2540));
  orx  g2513(.a(n2540), .b(n857), .O(n2541));
  andx g2514(.a(n2541), .b(n278), .O(n2542));
  andx g2515(.a(n2165), .b(n1352), .O(n2543));
  orx  g2516(.a(n2543), .b(n2542), .O(n2544));
  andx g2517(.a(n1926), .b(n1006), .O(n2545));
  andx g2518(.a(n2545), .b(n1387), .O(n2546));
  andx g2519(.a(n2486), .b(n576), .O(n2547));
  orx  g2520(.a(n2547), .b(n2546), .O(n2548));
  orx  g2521(.a(n2548), .b(n2544), .O(n2549));
  orx  g2522(.a(n2549), .b(n2539), .O(n2550));
  orx  g2523(.a(n2550), .b(n2532), .O(n2551));
  andx g2524(.a(n2510), .b(n858), .O(n2552));
  orx  g2525(.a(n178), .b(n139), .O(n2553));
  andx g2526(.a(n2553), .b(n1610), .O(n2554));
  orx  g2527(.a(n2554), .b(n2552), .O(n2555));
  andx g2528(.a(n1355), .b(n312), .O(n2556));
  andx g2529(.a(n920), .b(n267), .O(n2557));
  orx  g2530(.a(n2557), .b(n2556), .O(n2558));
  orx  g2531(.a(n2558), .b(n2555), .O(n2559));
  andx g2532(.a(n534), .b(n109), .O(n2560));
  andx g2533(.a(n2560), .b(n958), .O(n2561));
  andx g2534(.a(n1825), .b(n33), .O(n2562));
  orx  g2535(.a(n2562), .b(n2561), .O(n2563));
  andx g2536(.a(n397), .b(n37), .O(n2564));
  andx g2537(.a(n2564), .b(n146), .O(n2565));
  andx g2538(.a(n2565), .b(n701), .O(n2566));
  andx g2539(.a(n2560), .b(n956), .O(n2567));
  orx  g2540(.a(n2567), .b(n2566), .O(n2568));
  orx  g2541(.a(n2568), .b(n2563), .O(n2569));
  orx  g2542(.a(n2569), .b(n2559), .O(n2570));
  andx g2543(.a(n2540), .b(n859), .O(n2571));
  andx g2544(.a(n2485), .b(n1062), .O(n2572));
  orx  g2545(.a(n2572), .b(n2571), .O(n2573));
  orx  g2546(.a(n2573), .b(n572), .O(n2574));
  andx g2547(.a(n957), .b(n59), .O(n2575));
  andx g2548(.a(n2575), .b(n2510), .O(n2576));
  andx g2549(.a(n2515), .b(n107), .O(n2577));
  orx  g2550(.a(n2577), .b(n2576), .O(n2578));
  andx g2551(.a(n2471), .b(n33), .O(n2579));
  orx  g2552(.a(n2579), .b(n2426), .O(n2580));
  orx  g2553(.a(n2580), .b(n2578), .O(n2581));
  orx  g2554(.a(n2581), .b(n2574), .O(n2582));
  orx  g2555(.a(n2582), .b(n2570), .O(n2583));
  andx g2556(.a(n1926), .b(n110), .O(n2584));
  andx g2557(.a(n2584), .b(n582), .O(n2585));
  orx  g2558(.a(n2585), .b(n2457), .O(n2586));
  orx  g2559(.a(n2166), .b(n2088), .O(n2587));
  orx  g2560(.a(n2587), .b(n2586), .O(n2588));
  andx g2561(.a(n2471), .b(n123), .O(n2589));
  andx g2562(.a(n914), .b(n808), .O(n2590));
  orx  g2563(.a(n2590), .b(n2589), .O(n2591));
  andx g2564(.a(n2470), .b(n1825), .O(n2592));
  orx  g2565(.a(n2592), .b(n913), .O(n2593));
  orx  g2566(.a(n2593), .b(n2591), .O(n2594));
  orx  g2567(.a(n2594), .b(n2588), .O(n2595));
  andx g2568(.a(n2275), .b(n1062), .O(n2596));
  orx  g2569(.a(n2596), .b(n851), .O(n2597));
  andx g2570(.a(n2519), .b(n932), .O(n2598));
  orx  g2571(.a(n2598), .b(n2283), .O(n2599));
  orx  g2572(.a(n2599), .b(n2597), .O(n2600));
  andx g2573(.a(n1610), .b(n940), .O(n2601));
  andx g2574(.a(n2584), .b(n914), .O(n2602));
  orx  g2575(.a(n2602), .b(n2601), .O(n2603));
  andx g2576(.a(n2535), .b(n908), .O(n2604));
  andx g2577(.a(n2500), .b(n47), .O(n2605));
  orx  g2578(.a(n2605), .b(n2604), .O(n2606));
  orx  g2579(.a(n2606), .b(n2603), .O(n2607));
  orx  g2580(.a(n2607), .b(n2600), .O(n2608));
  orx  g2581(.a(n2608), .b(n2595), .O(n2609));
  orx  g2582(.a(n2609), .b(n2583), .O(n2610));
  orx  g2583(.a(n2610), .b(n2551), .O(n2611));
  orx  g2584(.a(n2611), .b(n2508), .O(n2612));
  orx  g2585(.a(n2612), .b(n2479), .O(po11));
  andx g2586(.a(n213), .b(pi00), .O(n2614));
  andx g2587(.a(n2614), .b(n1234), .O(n2615));
  andx g2588(.a(n216), .b(n77), .O(n2616));
  andx g2589(.a(n2616), .b(n1962), .O(n2617));
  orx  g2590(.a(n2617), .b(n2615), .O(n2618));
  andx g2591(.a(n1968), .b(n804), .O(n2619));
  andx g2592(.a(n502), .b(n71), .O(n2620));
  andx g2593(.a(n2620), .b(n1925), .O(n2621));
  orx  g2594(.a(n2621), .b(n2619), .O(n2622));
  orx  g2595(.a(n2622), .b(n2618), .O(n2623));
  andx g2596(.a(n100), .b(n77), .O(n2624));
  andx g2597(.a(n2624), .b(n82), .O(n2625));
  andx g2598(.a(n2625), .b(n858), .O(n2626));
  andx g2599(.a(n419), .b(n74), .O(n2627));
  andx g2600(.a(n2627), .b(n81), .O(n2628));
  andx g2601(.a(pi07), .b(n37), .O(n2629));
  andx g2602(.a(n2629), .b(n36), .O(n2630));
  andx g2603(.a(n2630), .b(n2628), .O(n2631));
  orx  g2604(.a(n2631), .b(n2626), .O(n2632));
  andx g2605(.a(n198), .b(n36), .O(n2633));
  andx g2606(.a(n81), .b(n48), .O(n2634));
  andx g2607(.a(n2634), .b(pi09), .O(n2635));
  orx  g2608(.a(n2635), .b(n2633), .O(n2636));
  andx g2609(.a(n2636), .b(n1481), .O(n2637));
  orx  g2610(.a(pi09), .b(pi08), .O(n2638));
  invx g2611(.a(n2638), .O(n2639));
  andx g2612(.a(n2639), .b(pi07), .O(n2640));
  andx g2613(.a(n2640), .b(n872), .O(n2641));
  andx g2614(.a(n2641), .b(n177), .O(n2642));
  orx  g2615(.a(n2642), .b(n2637), .O(n2643));
  orx  g2616(.a(n2643), .b(n2632), .O(n2644));
  orx  g2617(.a(n2644), .b(n2623), .O(n2645));
  andx g2618(.a(n1523), .b(n310), .O(n2646));
  andx g2619(.a(n108), .b(n563), .O(n2647));
  andx g2620(.a(n2371), .b(n1898), .O(n2648));
  andx g2621(.a(n2648), .b(n2647), .O(n2649));
  andx g2622(.a(pi08), .b(n41), .O(n2650));
  andx g2623(.a(n2650), .b(pi01), .O(n2651));
  andx g2624(.a(n2651), .b(n2625), .O(n2652));
  orx  g2625(.a(n2652), .b(n2649), .O(n2653));
  orx  g2626(.a(n2653), .b(n2646), .O(n2654));
  andx g2627(.a(n1962), .b(n104), .O(n2655));
  andx g2628(.a(n100), .b(n72), .O(n2656));
  andx g2629(.a(n2656), .b(n1925), .O(n2657));
  orx  g2630(.a(n2657), .b(n2655), .O(n2658));
  andx g2631(.a(n297), .b(n90), .O(n2659));
  andx g2632(.a(n2659), .b(n755), .O(n2660));
  andx g2633(.a(n100), .b(n563), .O(n2661));
  andx g2634(.a(n2661), .b(n2629), .O(n2662));
  andx g2635(.a(n2662), .b(n1899), .O(n2663));
  orx  g2636(.a(n2663), .b(n2660), .O(n2664));
  orx  g2637(.a(n2664), .b(n2658), .O(n2665));
  orx  g2638(.a(n2665), .b(n2654), .O(n2666));
  orx  g2639(.a(n2666), .b(n2645), .O(n2667));
  andx g2640(.a(n1952), .b(pi00), .O(n2668));
  andx g2641(.a(n60), .b(n48), .O(n2669));
  andx g2642(.a(n2669), .b(n2668), .O(n2670));
  andx g2643(.a(n2670), .b(n31), .O(n2671));
  andx g2644(.a(n910), .b(n85), .O(n2672));
  andx g2645(.a(n2672), .b(n771), .O(n2673));
  orx  g2646(.a(n2673), .b(n2671), .O(n2674));
  andx g2647(.a(n755), .b(n242), .O(n2675));
  andx g2648(.a(n2675), .b(n300), .O(n2676));
  andx g2649(.a(n82), .b(n74), .O(n2677));
  andx g2650(.a(n2677), .b(pi08), .O(n2678));
  andx g2651(.a(n2678), .b(n181), .O(n2679));
  orx  g2652(.a(n2679), .b(n2676), .O(n2680));
  orx  g2653(.a(n2680), .b(n2674), .O(n2681));
  andx g2654(.a(n73), .b(pi08), .O(n2682));
  andx g2655(.a(n2682), .b(n29), .O(n2683));
  andx g2656(.a(n2683), .b(n2227), .O(n2684));
  andx g2657(.a(n910), .b(n28), .O(n2685));
  orx  g2658(.a(n2685), .b(n386), .O(n2686));
  andx g2659(.a(n2686), .b(n30), .O(n2687));
  orx  g2660(.a(n2687), .b(n2684), .O(n2688));
  andx g2661(.a(n580), .b(pi07), .O(n2689));
  andx g2662(.a(n2689), .b(n879), .O(n2690));
  andx g2663(.a(n2690), .b(n596), .O(n2691));
  andx g2664(.a(n992), .b(n109), .O(n2692));
  orx  g2665(.a(n2692), .b(n2691), .O(n2693));
  orx  g2666(.a(n2693), .b(n2688), .O(n2694));
  orx  g2667(.a(n2694), .b(n2681), .O(n2695));
  andx g2668(.a(n502), .b(n397), .O(n2696));
  orx  g2669(.a(n48), .b(pi04), .O(n2697));
  andx g2670(.a(n2697), .b(pi01), .O(n2698));
  andx g2671(.a(n2698), .b(n2696), .O(n2699));
  andx g2672(.a(n108), .b(n36), .O(n2700));
  andx g2673(.a(n2700), .b(n2648), .O(n2701));
  orx  g2674(.a(n2701), .b(n2699), .O(n2702));
  andx g2675(.a(n48), .b(pi03), .O(n2703));
  andx g2676(.a(n2703), .b(n36), .O(n2704));
  orx  g2677(.a(n99), .b(pi09), .O(n2705));
  andx g2678(.a(n2705), .b(n74), .O(n2706));
  andx g2679(.a(n2706), .b(n2096), .O(n2707));
  andx g2680(.a(n2707), .b(n2704), .O(n2708));
  andx g2681(.a(n2625), .b(n580), .O(n2709));
  orx  g2682(.a(n2709), .b(n2708), .O(n2710));
  orx  g2683(.a(n2710), .b(n2702), .O(n2711));
  andx g2684(.a(n1963), .b(n1194), .O(n2712));
  andx g2685(.a(n230), .b(n29), .O(n2713));
  andx g2686(.a(n2713), .b(n2712), .O(n2714));
  andx g2687(.a(n2670), .b(n266), .O(n2715));
  orx  g2688(.a(n2715), .b(n2714), .O(n2716));
  andx g2689(.a(n41), .b(n37), .O(n2717));
  andx g2690(.a(n2717), .b(pi02), .O(n2718));
  andx g2691(.a(n75), .b(pi06), .O(n2719));
  andx g2692(.a(n2719), .b(n2718), .O(n2720));
  andx g2693(.a(n2647), .b(n992), .O(n2721));
  orx  g2694(.a(n2721), .b(n2720), .O(n2722));
  orx  g2695(.a(n2722), .b(n2716), .O(n2723));
  orx  g2696(.a(n2723), .b(n2711), .O(n2724));
  orx  g2697(.a(n2724), .b(n2695), .O(n2725));
  andx g2698(.a(n100), .b(n28), .O(n2726));
  andx g2699(.a(n2726), .b(n1962), .O(n2727));
  andx g2700(.a(n301), .b(n71), .O(n2728));
  andx g2701(.a(n2682), .b(n81), .O(n2729));
  orx  g2702(.a(n2729), .b(n2728), .O(n2730));
  orx  g2703(.a(n41), .b(n59), .O(n2731));
  andx g2704(.a(n48), .b(n36), .O(n2732));
  andx g2705(.a(n2732), .b(n2731), .O(n2733));
  andx g2706(.a(n2733), .b(n29), .O(n2734));
  andx g2707(.a(n2734), .b(n2730), .O(n2735));
  orx  g2708(.a(n2735), .b(n2727), .O(n2736));
  andx g2709(.a(n74), .b(n71), .O(n2737));
  andx g2710(.a(n2737), .b(n1981), .O(n2738));
  andx g2711(.a(n2717), .b(n620), .O(n2739));
  andx g2712(.a(n2739), .b(n515), .O(n2740));
  orx  g2713(.a(n2740), .b(n2738), .O(n2741));
  orx  g2714(.a(n2741), .b(n2736), .O(n2742));
  andx g2715(.a(n2627), .b(pi10), .O(n2743));
  andx g2716(.a(n2743), .b(n2718), .O(n2744));
  andx g2717(.a(n216), .b(n99), .O(n2745));
  andx g2718(.a(n2745), .b(n1962), .O(n2746));
  orx  g2719(.a(n2746), .b(n2744), .O(n2747));
  andx g2720(.a(n59), .b(n36), .O(n2748));
  andx g2721(.a(n2748), .b(pi07), .O(n2749));
  orx  g2722(.a(n2749), .b(n2124), .O(n2750));
  andx g2723(.a(n2750), .b(n2737), .O(n2751));
  andx g2724(.a(n1968), .b(n119), .O(n2752));
  orx  g2725(.a(n2752), .b(n2751), .O(n2753));
  orx  g2726(.a(n2753), .b(n2747), .O(n2754));
  orx  g2727(.a(n2754), .b(n2742), .O(n2755));
  andx g2728(.a(n100), .b(n71), .O(n2756));
  andx g2729(.a(n2756), .b(n28), .O(n2757));
  andx g2730(.a(n2757), .b(n1925), .O(n2758));
  andx g2731(.a(n2656), .b(n1962), .O(n2759));
  orx  g2732(.a(n2759), .b(n2758), .O(n2760));
  andx g2733(.a(n583), .b(n74), .O(n2761));
  andx g2734(.a(pi06), .b(n59), .O(n2762));
  andx g2735(.a(n2762), .b(n36), .O(n2763));
  orx  g2736(.a(n2763), .b(n2718), .O(n2764));
  andx g2737(.a(n2764), .b(n2761), .O(n2765));
  andx g2738(.a(n277), .b(n229), .O(n2766));
  andx g2739(.a(n2766), .b(n2712), .O(n2767));
  orx  g2740(.a(n2767), .b(n2765), .O(n2768));
  orx  g2741(.a(n2768), .b(n2760), .O(n2769));
  andx g2742(.a(n2641), .b(n1331), .O(n2770));
  andx g2743(.a(n108), .b(pi00), .O(n2771));
  andx g2744(.a(n2771), .b(n2648), .O(n2772));
  orx  g2745(.a(n2772), .b(n2770), .O(n2773));
  andx g2746(.a(n28), .b(n77), .O(n2774));
  orx  g2747(.a(n2774), .b(n120), .O(n2775));
  andx g2748(.a(n2775), .b(n100), .O(n2776));
  andx g2749(.a(n2776), .b(n591), .O(n2777));
  andx g2750(.a(n2700), .b(n992), .O(n2778));
  orx  g2751(.a(n2778), .b(n2777), .O(n2779));
  orx  g2752(.a(n2779), .b(n2773), .O(n2780));
  orx  g2753(.a(n2780), .b(n2769), .O(n2781));
  orx  g2754(.a(n2781), .b(n2755), .O(n2782));
  orx  g2755(.a(n2782), .b(n2725), .O(n2783));
  orx  g2756(.a(n2783), .b(n2667), .O(n2784));
  andx g2757(.a(n910), .b(n100), .O(n2785));
  andx g2758(.a(n2785), .b(n385), .O(n2786));
  andx g2759(.a(n2732), .b(pi09), .O(n2787));
  andx g2760(.a(n2787), .b(n162), .O(n2788));
  orx  g2761(.a(n2788), .b(n2786), .O(n2789));
  andx g2762(.a(pi08), .b(n59), .O(n2790));
  andx g2763(.a(n2790), .b(n36), .O(n2791));
  andx g2764(.a(n2791), .b(n297), .O(n2792));
  andx g2765(.a(n397), .b(n36), .O(n2793));
  andx g2766(.a(n2793), .b(n502), .O(n2794));
  orx  g2767(.a(n2794), .b(n2792), .O(n2795));
  orx  g2768(.a(n2795), .b(n2789), .O(n2796));
  andx g2769(.a(n1197), .b(pi05), .O(n2797));
  andx g2770(.a(n2797), .b(n103), .O(n2798));
  andx g2771(.a(n1905), .b(n2697), .O(n2799));
  andx g2772(.a(n2799), .b(n2661), .O(n2800));
  orx  g2773(.a(n2800), .b(n2798), .O(n2801));
  andx g2774(.a(n2624), .b(n134), .O(n2802));
  andx g2775(.a(n30), .b(n77), .O(n2803));
  andx g2776(.a(n2803), .b(n2019), .O(n2804));
  orx  g2777(.a(n2804), .b(n2802), .O(n2805));
  orx  g2778(.a(n2805), .b(n2801), .O(n2806));
  orx  g2779(.a(n2806), .b(n2796), .O(n2807));
  andx g2780(.a(n2718), .b(n297), .O(n2808));
  andx g2781(.a(n2803), .b(n2133), .O(n2809));
  orx  g2782(.a(n2809), .b(n2808), .O(n2810));
  andx g2783(.a(n134), .b(n101), .O(n2811));
  andx g2784(.a(n74), .b(n48), .O(n2812));
  andx g2785(.a(n2812), .b(n2633), .O(n2813));
  orx  g2786(.a(n2813), .b(n2811), .O(n2814));
  orx  g2787(.a(n2814), .b(n2810), .O(n2815));
  andx g2788(.a(n133), .b(pi09), .O(n2816));
  andx g2789(.a(n2816), .b(n162), .O(n2817));
  andx g2790(.a(n2717), .b(n59), .O(n2818));
  andx g2791(.a(n2818), .b(n119), .O(n2819));
  orx  g2792(.a(n2819), .b(n2817), .O(n2820));
  andx g2793(.a(n100), .b(pi06), .O(n2821));
  andx g2794(.a(n2821), .b(n1953), .O(n2822));
  andx g2795(.a(n2717), .b(n276), .O(n2823));
  andx g2796(.a(n2823), .b(n119), .O(n2824));
  orx  g2797(.a(n2824), .b(n2822), .O(n2825));
  orx  g2798(.a(n2825), .b(n2820), .O(n2826));
  orx  g2799(.a(n2826), .b(n2815), .O(n2827));
  orx  g2800(.a(n2827), .b(n2807), .O(n2828));
  andx g2801(.a(n29), .b(n71), .O(n2829));
  andx g2802(.a(n2829), .b(n113), .O(n2830));
  andx g2803(.a(n213), .b(pi02), .O(n2831));
  andx g2804(.a(n2831), .b(n2830), .O(n2832));
  andx g2805(.a(n2748), .b(n74), .O(n2833));
  andx g2806(.a(n2833), .b(n420), .O(n2834));
  orx  g2807(.a(n2834), .b(n2832), .O(n2835));
  andx g2808(.a(n385), .b(n74), .O(n2836));
  andx g2809(.a(n2836), .b(n2718), .O(n2837));
  orx  g2810(.a(n59), .b(n36), .O(n2838));
  andx g2811(.a(n1197), .b(n100), .O(n2839));
  andx g2812(.a(n2839), .b(n2838), .O(n2840));
  orx  g2813(.a(n2840), .b(n2837), .O(n2841));
  orx  g2814(.a(n2841), .b(n2835), .O(n2842));
  andx g2815(.a(n315), .b(n242), .O(n2843));
  andx g2816(.a(pi09), .b(n48), .O(n2844));
  andx g2817(.a(n2829), .b(n479), .O(n2845));
  andx g2818(.a(n2845), .b(n2844), .O(n2846));
  orx  g2819(.a(n2846), .b(n2843), .O(n2847));
  andx g2820(.a(n2096), .b(n30), .O(n2848));
  andx g2821(.a(n49), .b(n276), .O(n2849));
  andx g2822(.a(n2849), .b(n2848), .O(n2850));
  andx g2823(.a(n385), .b(n30), .O(n2851));
  andx g2824(.a(n2851), .b(n563), .O(n2852));
  orx  g2825(.a(n2852), .b(n2850), .O(n2853));
  orx  g2826(.a(n2853), .b(n2847), .O(n2854));
  orx  g2827(.a(n2854), .b(n2842), .O(n2855));
  andx g2828(.a(n2818), .b(n2371), .O(n2856));
  andx g2829(.a(n1197), .b(n41), .O(n2857));
  andx g2830(.a(n2857), .b(n101), .O(n2858));
  orx  g2831(.a(n2858), .b(n2856), .O(n2859));
  andx g2832(.a(n99), .b(n37), .O(n2860));
  andx g2833(.a(n2860), .b(n2839), .O(n2861));
  andx g2834(.a(n1197), .b(n74), .O(n2862));
  andx g2835(.a(n2862), .b(n147), .O(n2863));
  orx  g2836(.a(n2863), .b(n2861), .O(n2864));
  orx  g2837(.a(n2864), .b(n2859), .O(n2865));
  andx g2838(.a(n1952), .b(pi02), .O(n2866));
  andx g2839(.a(n73), .b(n41), .O(n2867));
  andx g2840(.a(n2867), .b(n2829), .O(n2868));
  andx g2841(.a(n2868), .b(n2866), .O(n2869));
  andx g2842(.a(n2627), .b(n1953), .O(n2870));
  orx  g2843(.a(n2870), .b(n2869), .O(n2871));
  andx g2844(.a(n2729), .b(n401), .O(n2872));
  andx g2845(.a(n2797), .b(n596), .O(n2873));
  orx  g2846(.a(n2873), .b(n2872), .O(n2874));
  orx  g2847(.a(n2874), .b(n2871), .O(n2875));
  orx  g2848(.a(n2875), .b(n2865), .O(n2876));
  orx  g2849(.a(n2876), .b(n2855), .O(n2877));
  orx  g2850(.a(n2877), .b(n2828), .O(n2878));
  andx g2851(.a(n2634), .b(n119), .O(n2879));
  andx g2852(.a(n100), .b(n48), .O(n2880));
  andx g2853(.a(n2717), .b(n2838), .O(n2881));
  andx g2854(.a(n2881), .b(n2880), .O(n2882));
  orx  g2855(.a(n2882), .b(n2879), .O(n2883));
  andx g2856(.a(n1908), .b(n1006), .O(n2884));
  andx g2857(.a(n2851), .b(n2614), .O(n2885));
  orx  g2858(.a(n2885), .b(n2884), .O(n2886));
  orx  g2859(.a(n2886), .b(n2883), .O(n2887));
  andx g2860(.a(n253), .b(n30), .O(n2888));
  andx g2861(.a(n2888), .b(n591), .O(n2889));
  andx g2862(.a(n29), .b(n48), .O(n2890));
  andx g2863(.a(n2890), .b(n51), .O(n2891));
  orx  g2864(.a(n41), .b(pi03), .O(n2892));
  andx g2865(.a(n37), .b(n276), .O(n2893));
  andx g2866(.a(n2893), .b(n2892), .O(n2894));
  andx g2867(.a(n2894), .b(n2891), .O(n2895));
  orx  g2868(.a(n2895), .b(n2889), .O(n2896));
  andx g2869(.a(n2726), .b(n1197), .O(n2897));
  andx g2870(.a(n2763), .b(n297), .O(n2898));
  orx  g2871(.a(n2898), .b(n2897), .O(n2899));
  orx  g2872(.a(n2899), .b(n2896), .O(n2900));
  orx  g2873(.a(n2900), .b(n2887), .O(n2901));
  andx g2874(.a(n2677), .b(n386), .O(n2902));
  andx g2875(.a(n1898), .b(n74), .O(n2903));
  andx g2876(.a(n2903), .b(n942), .O(n2904));
  orx  g2877(.a(n2904), .b(n2902), .O(n2905));
  andx g2878(.a(n28), .b(n48), .O(n2906));
  andx g2879(.a(n2906), .b(n30), .O(n2907));
  andx g2880(.a(n2907), .b(n2818), .O(n2908));
  orx  g2881(.a(n48), .b(pi05), .O(n2909));
  andx g2882(.a(n253), .b(n2909), .O(n2910));
  andx g2883(.a(n2910), .b(n2862), .O(n2911));
  orx  g2884(.a(n2911), .b(n2908), .O(n2912));
  orx  g2885(.a(n2912), .b(n2905), .O(n2913));
  andx g2886(.a(n2862), .b(n177), .O(n2914));
  andx g2887(.a(n2891), .b(n2818), .O(n2915));
  orx  g2888(.a(n2915), .b(n2914), .O(n2916));
  andx g2889(.a(n2677), .b(n2124), .O(n2917));
  andx g2890(.a(n30), .b(n41), .O(n2918));
  andx g2891(.a(n2638), .b(n385), .O(n2919));
  andx g2892(.a(n2919), .b(n2918), .O(n2920));
  orx  g2893(.a(n2920), .b(n2917), .O(n2921));
  orx  g2894(.a(n2921), .b(n2916), .O(n2922));
  orx  g2895(.a(n2922), .b(n2913), .O(n2923));
  orx  g2896(.a(n2923), .b(n2901), .O(n2924));
  andx g2897(.a(n2888), .b(n2849), .O(n2925));
  andx g2898(.a(n133), .b(n563), .O(n2926));
  andx g2899(.a(n2926), .b(n103), .O(n2927));
  orx  g2900(.a(n2927), .b(n2925), .O(n2928));
  andx g2901(.a(n591), .b(n101), .O(n2929));
  andx g2902(.a(n770), .b(n563), .O(n2930));
  andx g2903(.a(n2930), .b(n2756), .O(n2931));
  orx  g2904(.a(n2931), .b(n2929), .O(n2932));
  orx  g2905(.a(n2932), .b(n2928), .O(n2933));
  andx g2906(.a(n28), .b(pi05), .O(n2934));
  andx g2907(.a(n2934), .b(n74), .O(n2935));
  andx g2908(.a(n2935), .b(n1953), .O(n2936));
  andx g2909(.a(n2844), .b(pi00), .O(n2937));
  andx g2910(.a(n2937), .b(n162), .O(n2938));
  orx  g2911(.a(n2938), .b(n2936), .O(n2939));
  andx g2912(.a(n133), .b(n36), .O(n2940));
  andx g2913(.a(n2940), .b(n2627), .O(n2941));
  andx g2914(.a(n2890), .b(n2682), .O(n2942));
  andx g2915(.a(n2942), .b(n2718), .O(n2943));
  orx  g2916(.a(n2943), .b(n2941), .O(n2944));
  orx  g2917(.a(n2944), .b(n2939), .O(n2945));
  orx  g2918(.a(n2945), .b(n2933), .O(n2946));
  andx g2919(.a(n2823), .b(n131), .O(n2947));
  orx  g2920(.a(pi04), .b(n59), .O(n2948));
  andx g2921(.a(n2844), .b(n2948), .O(n2949));
  andx g2922(.a(n2949), .b(n162), .O(n2950));
  orx  g2923(.a(n2950), .b(n2947), .O(n2951));
  andx g2924(.a(n180), .b(n36), .O(n2952));
  andx g2925(.a(n2952), .b(n2830), .O(n2953));
  andx g2926(.a(n590), .b(n36), .O(n2954));
  andx g2927(.a(n2954), .b(n1836), .O(n2955));
  orx  g2928(.a(n2955), .b(n2953), .O(n2956));
  orx  g2929(.a(n2956), .b(n2951), .O(n2957));
  andx g2930(.a(n2844), .b(n74), .O(n2958));
  andx g2931(.a(n2958), .b(n2718), .O(n2959));
  andx g2932(.a(n438), .b(n100), .O(n2960));
  andx g2933(.a(n2960), .b(n1935), .O(n2961));
  orx  g2934(.a(n2961), .b(n2959), .O(n2962));
  orx  g2935(.a(n81), .b(pi09), .O(n2963));
  andx g2936(.a(n2963), .b(n30), .O(n2964));
  andx g2937(.a(n2964), .b(n2818), .O(n2965));
  andx g2938(.a(n2918), .b(n1953), .O(n2966));
  orx  g2939(.a(n2966), .b(n2965), .O(n2967));
  orx  g2940(.a(n2967), .b(n2962), .O(n2968));
  orx  g2941(.a(n2968), .b(n2957), .O(n2969));
  orx  g2942(.a(n2969), .b(n2946), .O(n2970));
  orx  g2943(.a(n2970), .b(n2924), .O(n2971));
  orx  g2944(.a(n2971), .b(n2878), .O(n2972));
  andx g2945(.a(n2954), .b(n2743), .O(n2973));
  andx g2946(.a(n2903), .b(pi07), .O(n2974));
  andx g2947(.a(n2974), .b(n64), .O(n2975));
  orx  g2948(.a(n2975), .b(n2973), .O(n2976));
  orx  g2949(.a(n2954), .b(n2940), .O(n2977));
  andx g2950(.a(n297), .b(pi08), .O(n2978));
  andx g2951(.a(n2978), .b(n2977), .O(n2979));
  andx g2952(.a(pi07), .b(pi02), .O(n2980));
  andx g2953(.a(n2980), .b(n1008), .O(n2981));
  orx  g2954(.a(n2981), .b(n2700), .O(n2982));
  andx g2955(.a(n2982), .b(n2672), .O(n2983));
  orx  g2956(.a(n2983), .b(n2979), .O(n2984));
  orx  g2957(.a(n2984), .b(n2976), .O(n2985));
  andx g2958(.a(n2650), .b(n85), .O(n2986));
  andx g2959(.a(n2986), .b(n2866), .O(n2987));
  andx g2960(.a(pi10), .b(n71), .O(n2988));
  andx g2961(.a(n2988), .b(n74), .O(n2989));
  andx g2962(.a(n2989), .b(n48), .O(n2990));
  andx g2963(.a(n2990), .b(n2718), .O(n2991));
  orx  g2964(.a(n2991), .b(n2987), .O(n2992));
  orx  g2965(.a(n41), .b(n37), .O(n2993));
  orx  g2966(.a(n2993), .b(n28), .O(n2994));
  andx g2967(.a(n2994), .b(n910), .O(n2995));
  andx g2968(.a(n2995), .b(n2624), .O(n2996));
  orx  g2969(.a(n2844), .b(n187), .O(n2997));
  andx g2970(.a(n2997), .b(n2625), .O(n2998));
  orx  g2971(.a(n2998), .b(n2996), .O(n2999));
  orx  g2972(.a(n2999), .b(n2992), .O(n3000));
  orx  g2973(.a(n3000), .b(n2985), .O(n3001));
  orx  g2974(.a(n1288), .b(n109), .O(n3002));
  andx g2975(.a(n3002), .b(n1951), .O(n3003));
  orx  g2976(.a(n2907), .b(n2891), .O(n3004));
  andx g2977(.a(n3004), .b(n1968), .O(n3005));
  orx  g2978(.a(n3005), .b(n3003), .O(n3006));
  orx  g2979(.a(pi05), .b(n59), .O(n3007));
  andx g2980(.a(n3007), .b(n2696), .O(n3008));
  andx g2981(.a(n2762), .b(n1309), .O(n3009));
  andx g2982(.a(n3009), .b(n2712), .O(n3010));
  orx  g2983(.a(n3010), .b(n3008), .O(n3011));
  orx  g2984(.a(n3011), .b(n3006), .O(n3012));
  andx g2985(.a(n2717), .b(pi01), .O(n3013));
  orx  g2986(.a(n3013), .b(n591), .O(n3014));
  andx g2987(.a(n3014), .b(n2880), .O(n3015));
  andx g2988(.a(n2791), .b(n2743), .O(n3016));
  orx  g2989(.a(n3016), .b(n3015), .O(n3017));
  orx  g2990(.a(n2756), .b(n31), .O(n3018));
  andx g2991(.a(n3018), .b(n385), .O(n3019));
  andx g2992(.a(n1915), .b(n108), .O(n3020));
  andx g2993(.a(n3020), .b(n2648), .O(n3021));
  orx  g2994(.a(n3021), .b(n3019), .O(n3022));
  orx  g2995(.a(n3022), .b(n3017), .O(n3023));
  orx  g2996(.a(n3023), .b(n3012), .O(n3024));
  orx  g2997(.a(n3024), .b(n3001), .O(n3025));
  orx  g2998(.a(n2954), .b(n2718), .O(n3026));
  andx g2999(.a(n420), .b(n74), .O(n3027));
  andx g3000(.a(n3027), .b(n3026), .O(n3028));
  andx g3001(.a(n563), .b(n276), .O(n3029));
  andx g3002(.a(n3029), .b(n30), .O(n3030));
  andx g3003(.a(n36), .b(n563), .O(n3031));
  andx g3004(.a(n3031), .b(n100), .O(n3032));
  orx  g3005(.a(n3032), .b(n2851), .O(n3033));
  orx  g3006(.a(n3033), .b(n3030), .O(n3034));
  orx  g3007(.a(n3034), .b(n3028), .O(n3035));
  andx g3008(.a(n180), .b(n59), .O(n3036));
  orx  g3009(.a(n3036), .b(n2831), .O(n3037));
  andx g3010(.a(n3037), .b(n2678), .O(n3038));
  orx  g3011(.a(pi04), .b(pi03), .O(n3039));
  andx g3012(.a(n3039), .b(n213), .O(n3040));
  andx g3013(.a(n3040), .b(n1234), .O(n3041));
  orx  g3014(.a(n3041), .b(n3038), .O(n3042));
  orx  g3015(.a(n3042), .b(n3035), .O(n3043));
  andx g3016(.a(n2818), .b(n131), .O(n3044));
  andx g3017(.a(n73), .b(n71), .O(n3045));
  andx g3018(.a(n3045), .b(n1309), .O(n3046));
  andx g3019(.a(n3046), .b(n1953), .O(n3047));
  orx  g3020(.a(n3047), .b(n3044), .O(n3048));
  andx g3021(.a(n3036), .b(n2868), .O(n3049));
  andx g3022(.a(n3045), .b(n771), .O(n3050));
  orx  g3023(.a(n3050), .b(n3049), .O(n3051));
  orx  g3024(.a(n3051), .b(n3048), .O(n3052));
  andx g3025(.a(n133), .b(n73), .O(n3053));
  andx g3026(.a(n3053), .b(n253), .O(n3054));
  andx g3027(.a(n2989), .b(n2733), .O(n3055));
  orx  g3028(.a(n3055), .b(n3054), .O(n3056));
  andx g3029(.a(n216), .b(n134), .O(n3057));
  andx g3030(.a(n2737), .b(n386), .O(n3058));
  orx  g3031(.a(n3058), .b(n3057), .O(n3059));
  orx  g3032(.a(n3059), .b(n3056), .O(n3060));
  orx  g3033(.a(n3060), .b(n3052), .O(n3061));
  orx  g3034(.a(n3061), .b(n3043), .O(n3062));
  orx  g3035(.a(pi03), .b(n36), .O(n3063));
  andx g3036(.a(n2893), .b(n3063), .O(n3064));
  orx  g3037(.a(n3064), .b(n2668), .O(n3065));
  andx g3038(.a(n3065), .b(n2918), .O(n3066));
  andx g3039(.a(n2739), .b(n101), .O(n3067));
  orx  g3040(.a(n3067), .b(n3066), .O(n3068));
  andx g3041(.a(n2974), .b(n2704), .O(n3069));
  orx  g3042(.a(n1331), .b(n39), .O(n3070));
  andx g3043(.a(n3070), .b(n2862), .O(n3071));
  orx  g3044(.a(n3071), .b(n3069), .O(n3072));
  orx  g3045(.a(n3072), .b(n3068), .O(n3073));
  orx  g3046(.a(pi07), .b(pi05), .O(n3074));
  orx  g3047(.a(n3074), .b(n36), .O(n3075));
  andx g3048(.a(n1197), .b(n29), .O(n3076));
  andx g3049(.a(n3076), .b(n272), .O(n3077));
  andx g3050(.a(n3077), .b(n3075), .O(n3078));
  andx g3051(.a(n770), .b(pi02), .O(n3079));
  andx g3052(.a(n2732), .b(n77), .O(n3080));
  orx  g3053(.a(n3080), .b(n3079), .O(n3081));
  andx g3054(.a(n2829), .b(n301), .O(n3082));
  andx g3055(.a(n3082), .b(n3081), .O(n3083));
  orx  g3056(.a(n3083), .b(n3078), .O(n3084));
  orx  g3057(.a(n2564), .b(n1926), .O(n3085));
  andx g3058(.a(n3085), .b(n2785), .O(n3086));
  orx  g3059(.a(n214), .b(n181), .O(n3087));
  andx g3060(.a(n3087), .b(n2620), .O(n3088));
  orx  g3061(.a(n3088), .b(n3086), .O(n3089));
  orx  g3062(.a(n3089), .b(n3084), .O(n3090));
  orx  g3063(.a(n3090), .b(n3073), .O(n3091));
  orx  g3064(.a(n3091), .b(n3062), .O(n3092));
  orx  g3065(.a(n3092), .b(n3025), .O(n3093));
  orx  g3066(.a(n3093), .b(n2972), .O(n3094));
  andx g3067(.a(n38), .b(n563), .O(n3095));
  orx  g3068(.a(n2696), .b(n2625), .O(n3096));
  andx g3069(.a(n3096), .b(n3095), .O(n3097));
  andx g3070(.a(n621), .b(n36), .O(n3098));
  andx g3071(.a(n3098), .b(n879), .O(n3099));
  andx g3072(.a(n2639), .b(n81), .O(n3100));
  andx g3073(.a(n2980), .b(pi05), .O(n3101));
  andx g3074(.a(n3101), .b(n3100), .O(n3102));
  orx  g3075(.a(n3102), .b(n3099), .O(n3103));
  andx g3076(.a(n3103), .b(n421), .O(n3104));
  invx g3077(.a(n1811), .O(n3105));
  andx g3078(.a(n30), .b(pi05), .O(n3106));
  andx g3079(.a(n3106), .b(n3105), .O(n3107));
  orx  g3080(.a(n3107), .b(n162), .O(n3108));
  andx g3081(.a(n3108), .b(n1968), .O(n3109));
  orx  g3082(.a(n3109), .b(n3104), .O(n3110));
  orx  g3083(.a(n3110), .b(n3097), .O(n3111));
  orx  g3084(.a(pi12), .b(n81), .O(n3112));
  orx  g3085(.a(n3112), .b(n28), .O(n3113));
  andx g3086(.a(n2756), .b(n3113), .O(n3114));
  orx  g3087(.a(n3114), .b(n452), .O(n3115));
  andx g3088(.a(n3115), .b(n591), .O(n3116));
  orx  g3089(.a(n3026), .b(n1906), .O(n3117));
  orx  g3090(.a(n120), .b(n32), .O(n3118));
  andx g3091(.a(n74), .b(pi06), .O(n3119));
  andx g3092(.a(n3119), .b(n3118), .O(n3120));
  andx g3093(.a(n3120), .b(n3117), .O(n3121));
  orx  g3094(.a(n3121), .b(n3116), .O(n3122));
  andx g3095(.a(n2730), .b(pi13), .O(n3123));
  andx g3096(.a(n3123), .b(n1962), .O(n3124));
  andx g3097(.a(n2980), .b(n1007), .O(n3125));
  orx  g3098(.a(n1633), .b(n97), .O(n3126));
  orx  g3099(.a(n3126), .b(n3125), .O(n3127));
  andx g3100(.a(n3127), .b(n2628), .O(n3128));
  orx  g3101(.a(n3128), .b(n3124), .O(n3129));
  orx  g3102(.a(n3129), .b(n3122), .O(n3130));
  orx  g3103(.a(n119), .b(n101), .O(n3131));
  orx  g3104(.a(n3131), .b(n297), .O(n3132));
  andx g3105(.a(n2096), .b(pi08), .O(n3133));
  andx g3106(.a(n3133), .b(n3132), .O(n3134));
  andx g3107(.a(n2849), .b(n194), .O(n3135));
  orx  g3108(.a(n99), .b(n81), .O(n3136));
  andx g3109(.a(n3136), .b(n60), .O(n3137));
  andx g3110(.a(n3137), .b(n2668), .O(n3138));
  orx  g3111(.a(n3138), .b(n3135), .O(n3139));
  andx g3112(.a(n3139), .b(n30), .O(n3140));
  orx  g3113(.a(n3140), .b(n3134), .O(n3141));
  invx g3114(.a(n63), .O(n3142));
  orx  g3115(.a(n1008), .b(n59), .O(n3143));
  orx  g3116(.a(n3143), .b(n3142), .O(n3144));
  andx g3117(.a(n3144), .b(n1811), .O(n3145));
  andx g3118(.a(n3145), .b(n1259), .O(n3146));
  orx  g3119(.a(n41), .b(n36), .O(n3147));
  andx g3120(.a(n180), .b(n3147), .O(n3148));
  orx  g3121(.a(n3148), .b(n386), .O(n3149));
  orx  g3122(.a(n3149), .b(n2124), .O(n3150));
  andx g3123(.a(n3150), .b(n1974), .O(n3151));
  orx  g3124(.a(n3151), .b(n3146), .O(n3152));
  orx  g3125(.a(n3152), .b(n3141), .O(n3153));
  orx  g3126(.a(n3153), .b(n3130), .O(n3154));
  orx  g3127(.a(n3154), .b(n3111), .O(n3155));
  andx g3128(.a(n1974), .b(n1926), .O(n3156));
  andx g3129(.a(n1898), .b(n100), .O(n3157));
  andx g3130(.a(n3157), .b(n942), .O(n3158));
  orx  g3131(.a(n3158), .b(n3156), .O(n3159));
  andx g3132(.a(n2785), .b(n1494), .O(n3160));
  andx g3133(.a(n2829), .b(n241), .O(n3161));
  andx g3134(.a(n3161), .b(n3148), .O(n3162));
  orx  g3135(.a(n3162), .b(n3160), .O(n3163));
  orx  g3136(.a(n3163), .b(n3159), .O(n3164));
  andx g3137(.a(n201), .b(n37), .O(n3165));
  andx g3138(.a(n3165), .b(n492), .O(n3166));
  andx g3139(.a(n1932), .b(n279), .O(n3167));
  orx  g3140(.a(n3167), .b(n3166), .O(n3168));
  andx g3141(.a(n3079), .b(n2989), .O(n3169));
  andx g3142(.a(n2954), .b(n75), .O(n3170));
  orx  g3143(.a(n3170), .b(n3169), .O(n3171));
  orx  g3144(.a(n3171), .b(n3168), .O(n3172));
  orx  g3145(.a(n3172), .b(n3164), .O(n3173));
  orx  g3146(.a(n2733), .b(n2636), .O(n3174));
  andx g3147(.a(n201), .b(n74), .O(n3175));
  andx g3148(.a(n3175), .b(n3174), .O(n3176));
  andx g3149(.a(n2848), .b(n1233), .O(n3177));
  orx  g3150(.a(pi08), .b(n77), .O(n3178));
  andx g3151(.a(n133), .b(n3178), .O(n3179));
  andx g3152(.a(n3179), .b(n2661), .O(n3180));
  orx  g3153(.a(n3180), .b(n3177), .O(n3181));
  andx g3154(.a(n2748), .b(n1008), .O(n3182));
  andx g3155(.a(n3182), .b(n2627), .O(n3183));
  andx g3156(.a(n151), .b(n74), .O(n3184));
  andx g3157(.a(n2748), .b(n2993), .O(n3185));
  andx g3158(.a(n3185), .b(n3184), .O(n3186));
  orx  g3159(.a(n3186), .b(n3183), .O(n3187));
  orx  g3160(.a(n3187), .b(n3181), .O(n3188));
  orx  g3161(.a(n3188), .b(n3176), .O(n3189));
  orx  g3162(.a(n3189), .b(n3173), .O(n3190));
  andx g3163(.a(n2907), .b(n2823), .O(n3191));
  andx g3164(.a(n2839), .b(n858), .O(n3192));
  orx  g3165(.a(n3192), .b(n3191), .O(n3193));
  andx g3166(.a(n2907), .b(n2849), .O(n3194));
  andx g3167(.a(n1898), .b(pi04), .O(n3195));
  andx g3168(.a(n3195), .b(n2656), .O(n3196));
  orx  g3169(.a(n3196), .b(n3194), .O(n3197));
  orx  g3170(.a(n3197), .b(n3193), .O(n3198));
  orx  g3171(.a(pi10), .b(pi09), .O(n3199));
  andx g3172(.a(n3199), .b(n100), .O(n3200));
  andx g3173(.a(n3200), .b(n134), .O(n3201));
  andx g3174(.a(n3161), .b(n2793), .O(n3202));
  orx  g3175(.a(n3202), .b(n3201), .O(n3203));
  andx g3176(.a(n2656), .b(n591), .O(n3204));
  andx g3177(.a(n3095), .b(n2839), .O(n3205));
  orx  g3178(.a(n3205), .b(n3204), .O(n3206));
  orx  g3179(.a(n3206), .b(n3203), .O(n3207));
  orx  g3180(.a(n3207), .b(n3198), .O(n3208));
  andx g3181(.a(n3157), .b(n685), .O(n3209));
  andx g3182(.a(n2903), .b(n1288), .O(n3210));
  orx  g3183(.a(n3210), .b(n3209), .O(n3211));
  andx g3184(.a(n2761), .b(n2633), .O(n3212));
  andx g3185(.a(n2926), .b(n101), .O(n3213));
  orx  g3186(.a(n3213), .b(n3212), .O(n3214));
  orx  g3187(.a(n3214), .b(n3211), .O(n3215));
  andx g3188(.a(n1197), .b(n130), .O(n3216));
  andx g3189(.a(n3216), .b(n1481), .O(n3217));
  andx g3190(.a(n2930), .b(n2785), .O(n3218));
  orx  g3191(.a(n3218), .b(n3217), .O(n3219));
  andx g3192(.a(n2816), .b(n2661), .O(n3220));
  andx g3193(.a(n2940), .b(n75), .O(n3221));
  orx  g3194(.a(n3221), .b(n3220), .O(n3222));
  orx  g3195(.a(n3222), .b(n3219), .O(n3223));
  orx  g3196(.a(n3223), .b(n3215), .O(n3224));
  orx  g3197(.a(n3224), .b(n3208), .O(n3225));
  orx  g3198(.a(n3225), .b(n3190), .O(n3226));
  orx  g3199(.a(n2963), .b(pi08), .O(n3227));
  andx g3200(.a(n2823), .b(n3227), .O(n3228));
  andx g3201(.a(n2849), .b(n99), .O(n3229));
  orx  g3202(.a(n3229), .b(n3228), .O(n3230));
  andx g3203(.a(n3230), .b(n30), .O(n3231));
  orx  g3204(.a(n2762), .b(n2703), .O(n3232));
  orx  g3205(.a(n3232), .b(n1009), .O(n3233));
  andx g3206(.a(n3233), .b(pi07), .O(n3234));
  andx g3207(.a(n3234), .b(n1951), .O(n3235));
  orx  g3208(.a(n3235), .b(n3231), .O(n3236));
  orx  g3209(.a(n3046), .b(n2935), .O(n3237));
  orx  g3210(.a(pi11), .b(pi10), .O(n3238));
  orx  g3211(.a(n3238), .b(n28), .O(n3239));
  andx g3212(.a(n3239), .b(pi06), .O(n3240));
  andx g3213(.a(n3240), .b(n90), .O(n3241));
  andx g3214(.a(n3241), .b(n3237), .O(n3242));
  orx  g3215(.a(n2625), .b(n2097), .O(n3243));
  andx g3216(.a(n3243), .b(n2838), .O(n3244));
  orx  g3217(.a(n3244), .b(n3242), .O(n3245));
  orx  g3218(.a(n3245), .b(n3236), .O(n3246));
  andx g3219(.a(n1309), .b(n51), .O(n3247));
  orx  g3220(.a(n3247), .b(n2845), .O(n3248));
  orx  g3221(.a(n3248), .b(n3107), .O(n3249));
  andx g3222(.a(n3249), .b(n2849), .O(n3250));
  orx  g3223(.a(pi09), .b(n77), .O(n3251));
  orx  g3224(.a(n1560), .b(pi07), .O(n3252));
  andx g3225(.a(n3252), .b(n3251), .O(n3253));
  orx  g3226(.a(n3253), .b(n32), .O(n3254));
  andx g3227(.a(n2739), .b(n100), .O(n3255));
  andx g3228(.a(n3255), .b(n3254), .O(n3256));
  orx  g3229(.a(n3256), .b(n3250), .O(n3257));
  orx  g3230(.a(n2966), .b(n2718), .O(n3258));
  andx g3231(.a(n3258), .b(n1481), .O(n3259));
  orx  g3232(.a(n3026), .b(n2763), .O(n3260));
  invx g3233(.a(n878), .O(n3261));
  orx  g3234(.a(pi09), .b(pi06), .O(n3262));
  andx g3235(.a(n3262), .b(n3261), .O(n3263));
  andx g3236(.a(n3263), .b(n3184), .O(n3264));
  andx g3237(.a(n3264), .b(n3260), .O(n3265));
  orx  g3238(.a(n3265), .b(n3259), .O(n3266));
  orx  g3239(.a(n3266), .b(n3257), .O(n3267));
  orx  g3240(.a(n3267), .b(n3246), .O(n3268));
  orx  g3241(.a(n3268), .b(n3226), .O(n3269));
  orx  g3242(.a(n3269), .b(n3155), .O(n3270));
  orx  g3243(.a(n3270), .b(n3094), .O(n3271));
  orx  g3244(.a(n3271), .b(n2784), .O(po12));
  andx g3245(.a(n1981), .b(n1951), .O(n3273));
  andx g3246(.a(n2640), .b(n1942), .O(n3274));
  andx g3247(.a(n1177), .b(n134), .O(n3275));
  andx g3248(.a(n3275), .b(n3274), .O(n3276));
  orx  g3249(.a(n3276), .b(n3273), .O(n3277));
  orx  g3250(.a(n2009), .b(n1947), .O(n3278));
  orx  g3251(.a(n3278), .b(n3277), .O(n3279));
  andx g3252(.a(n2818), .b(n1913), .O(n3280));
  andx g3253(.a(n3280), .b(n1198), .O(n3281));
  andx g3254(.a(n3281), .b(n1417), .O(n3282));
  orx  g3255(.a(n3282), .b(n1978), .O(n3283));
  orx  g3256(.a(n3283), .b(n3279), .O(n3284));
  andx g3257(.a(n3100), .b(n258), .O(n3285));
  andx g3258(.a(n3285), .b(n1901), .O(n3286));
  orx  g3259(.a(n3286), .b(n2004), .O(n3287));
  orx  g3260(.a(n1930), .b(n1910), .O(n3288));
  orx  g3261(.a(n3288), .b(n3287), .O(n3289));
  orx  g3262(.a(n3289), .b(n2100), .O(n3290));
  orx  g3263(.a(n3290), .b(n3284), .O(n3291));
  orx  g3264(.a(n2230), .b(n1922), .O(n3292));
  orx  g3265(.a(n3292), .b(n1904), .O(n3293));
  orx  g3266(.a(n3293), .b(n1972), .O(n3294));
  orx  g3267(.a(n3294), .b(n3291), .O(po13));
endmodule


