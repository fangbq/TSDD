// Benchmark "top" written by ABC on Sun Jan 26 11:08:06 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93,
    pi94, pi95;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31;
  wire n128, n129, n130, n131, n132, n133, n134, n135, n136, n138, n139,
    n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n499,
    n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n615, n616, n617, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n739, n740, n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190;
  invx  g0000(.a(pi00), .O(n128));
  andx  g0001(.a(pi01), .b(n128), .O(n129));
  invx  g0002(.a(pi01), .O(n130));
  andx  g0003(.a(n130), .b(pi00), .O(n131));
  orx   g0004(.a(n131), .b(n129), .O(n132));
  invx  g0005(.a(n132), .O(n133));
  andx  g0006(.a(n133), .b(pi02), .O(n134));
  invx  g0007(.a(pi02), .O(n135));
  andx  g0008(.a(n132), .b(n135), .O(n136));
  orx   g0009(.a(n136), .b(n134), .O(po00));
  invx  g0010(.a(pi04), .O(n138));
  orx   g0011(.a(n130), .b(n128), .O(n139));
  andx  g0012(.a(n139), .b(pi03), .O(n140));
  invx  g0013(.a(pi03), .O(n141));
  andx  g0014(.a(pi01), .b(pi00), .O(n142));
  andx  g0015(.a(n142), .b(n141), .O(n143));
  orx   g0016(.a(n143), .b(n140), .O(n144));
  andx  g0017(.a(n144), .b(n138), .O(n145));
  andx  g0018(.a(pi04), .b(n141), .O(n146));
  andx  g0019(.a(n146), .b(n139), .O(n147));
  andx  g0020(.a(n142), .b(pi04), .O(n148));
  andx  g0021(.a(n148), .b(pi03), .O(n149));
  orx   g0022(.a(n149), .b(n147), .O(n150));
  orx   g0023(.a(n150), .b(n145), .O(n151));
  andx  g0024(.a(n132), .b(pi02), .O(n152));
  orx   g0025(.a(n152), .b(n151), .O(n153));
  orx   g0026(.a(n142), .b(n141), .O(n154));
  orx   g0027(.a(n139), .b(pi03), .O(n155));
  andx  g0028(.a(n155), .b(n154), .O(n156));
  orx   g0029(.a(n156), .b(pi04), .O(n157));
  orx   g0030(.a(n138), .b(pi03), .O(n158));
  orx   g0031(.a(n158), .b(n142), .O(n159));
  orx   g0032(.a(n139), .b(n138), .O(n160));
  orx   g0033(.a(n160), .b(n141), .O(n161));
  andx  g0034(.a(n161), .b(n159), .O(n162));
  andx  g0035(.a(n162), .b(n157), .O(n163));
  invx  g0036(.a(n152), .O(n164));
  orx   g0037(.a(n164), .b(n163), .O(n165));
  andx  g0038(.a(n165), .b(n153), .O(n166));
  invx  g0039(.a(n166), .O(n167));
  andx  g0040(.a(n167), .b(pi05), .O(n168));
  invx  g0041(.a(pi05), .O(n169));
  andx  g0042(.a(n166), .b(n169), .O(n170));
  orx   g0043(.a(n170), .b(n168), .O(po01));
  invx  g0044(.a(pi06), .O(n172));
  andx  g0045(.a(pi07), .b(n172), .O(n173));
  invx  g0046(.a(pi07), .O(n174));
  andx  g0047(.a(n174), .b(pi06), .O(n175));
  orx   g0048(.a(n175), .b(n173), .O(n176));
  orx   g0049(.a(n142), .b(pi04), .O(n177));
  andx  g0050(.a(n177), .b(pi03), .O(n178));
  orx   g0051(.a(n178), .b(n148), .O(n179));
  andx  g0052(.a(n179), .b(n176), .O(n180));
  invx  g0053(.a(n180), .O(n181));
  orx   g0054(.a(n179), .b(n176), .O(n182));
  andx  g0055(.a(n182), .b(n181), .O(n183));
  andx  g0056(.a(n183), .b(pi08), .O(n184));
  invx  g0057(.a(pi08), .O(n185));
  invx  g0058(.a(n183), .O(n186));
  andx  g0059(.a(n186), .b(n185), .O(n187));
  orx   g0060(.a(n187), .b(n184), .O(n188));
  andx  g0061(.a(n152), .b(n151), .O(n189));
  andx  g0062(.a(n153), .b(pi05), .O(n190));
  orx   g0063(.a(n190), .b(n189), .O(n191));
  andx  g0064(.a(n191), .b(n188), .O(n192));
  invx  g0065(.a(n188), .O(n193));
  andx  g0066(.a(n164), .b(n163), .O(n194));
  orx   g0067(.a(n194), .b(n169), .O(n195));
  andx  g0068(.a(n195), .b(n165), .O(n196));
  andx  g0069(.a(n196), .b(n193), .O(n197));
  orx   g0070(.a(n197), .b(n192), .O(po02));
  invx  g0071(.a(pi09), .O(n199));
  andx  g0072(.a(pi10), .b(n199), .O(n200));
  invx  g0073(.a(pi10), .O(n201));
  andx  g0074(.a(n201), .b(pi09), .O(n202));
  orx   g0075(.a(n202), .b(n200), .O(n203));
  orx   g0076(.a(n179), .b(pi06), .O(n204));
  andx  g0077(.a(n204), .b(pi07), .O(n205));
  andx  g0078(.a(n179), .b(pi06), .O(n206));
  orx   g0079(.a(n206), .b(n205), .O(n207));
  andx  g0080(.a(n207), .b(n203), .O(n208));
  invx  g0081(.a(n208), .O(n209));
  orx   g0082(.a(n207), .b(n203), .O(n210));
  andx  g0083(.a(n210), .b(n209), .O(n211));
  andx  g0084(.a(n211), .b(pi11), .O(n212));
  invx  g0085(.a(pi11), .O(n213));
  invx  g0086(.a(n211), .O(n214));
  andx  g0087(.a(n214), .b(n213), .O(n215));
  orx   g0088(.a(n215), .b(n212), .O(n216));
  orx   g0089(.a(n191), .b(n183), .O(n217));
  andx  g0090(.a(n217), .b(pi08), .O(n218));
  andx  g0091(.a(n191), .b(n183), .O(n219));
  orx   g0092(.a(n219), .b(n218), .O(n220));
  andx  g0093(.a(n220), .b(n216), .O(n221));
  invx  g0094(.a(n216), .O(n222));
  andx  g0095(.a(n196), .b(n186), .O(n223));
  orx   g0096(.a(n223), .b(n185), .O(n224));
  orx   g0097(.a(n196), .b(n186), .O(n225));
  andx  g0098(.a(n225), .b(n224), .O(n226));
  andx  g0099(.a(n226), .b(n222), .O(n227));
  orx   g0100(.a(n227), .b(n221), .O(po03));
  invx  g0101(.a(pi12), .O(n229));
  andx  g0102(.a(pi13), .b(n229), .O(n230));
  invx  g0103(.a(pi13), .O(n231));
  andx  g0104(.a(n231), .b(pi12), .O(n232));
  orx   g0105(.a(n232), .b(n230), .O(n233));
  orx   g0106(.a(n207), .b(pi09), .O(n234));
  andx  g0107(.a(n234), .b(pi10), .O(n235));
  andx  g0108(.a(n207), .b(pi09), .O(n236));
  orx   g0109(.a(n236), .b(n235), .O(n237));
  andx  g0110(.a(n237), .b(n233), .O(n238));
  invx  g0111(.a(n238), .O(n239));
  orx   g0112(.a(n237), .b(n233), .O(n240));
  andx  g0113(.a(n240), .b(n239), .O(n241));
  andx  g0114(.a(n241), .b(pi14), .O(n242));
  invx  g0115(.a(pi14), .O(n243));
  invx  g0116(.a(n241), .O(n244));
  andx  g0117(.a(n244), .b(n243), .O(n245));
  orx   g0118(.a(n245), .b(n242), .O(n246));
  orx   g0119(.a(n220), .b(n211), .O(n247));
  andx  g0120(.a(n247), .b(pi11), .O(n248));
  andx  g0121(.a(n220), .b(n211), .O(n249));
  orx   g0122(.a(n249), .b(n248), .O(n250));
  andx  g0123(.a(n250), .b(n246), .O(n251));
  invx  g0124(.a(n246), .O(n252));
  andx  g0125(.a(n226), .b(n214), .O(n253));
  orx   g0126(.a(n253), .b(n213), .O(n254));
  orx   g0127(.a(n226), .b(n214), .O(n255));
  andx  g0128(.a(n255), .b(n254), .O(n256));
  andx  g0129(.a(n256), .b(n252), .O(n257));
  orx   g0130(.a(n257), .b(n251), .O(po04));
  invx  g0131(.a(pi15), .O(n259));
  andx  g0132(.a(pi16), .b(n259), .O(n260));
  invx  g0133(.a(pi16), .O(n261));
  andx  g0134(.a(n261), .b(pi15), .O(n262));
  orx   g0135(.a(n262), .b(n260), .O(n263));
  orx   g0136(.a(n237), .b(pi12), .O(n264));
  andx  g0137(.a(n264), .b(pi13), .O(n265));
  andx  g0138(.a(n237), .b(pi12), .O(n266));
  orx   g0139(.a(n266), .b(n265), .O(n267));
  andx  g0140(.a(n267), .b(n263), .O(n268));
  invx  g0141(.a(n268), .O(n269));
  orx   g0142(.a(n267), .b(n263), .O(n270));
  andx  g0143(.a(n270), .b(n269), .O(n271));
  andx  g0144(.a(n271), .b(pi17), .O(n272));
  invx  g0145(.a(pi17), .O(n273));
  invx  g0146(.a(n271), .O(n274));
  andx  g0147(.a(n274), .b(n273), .O(n275));
  orx   g0148(.a(n275), .b(n272), .O(n276));
  orx   g0149(.a(n250), .b(n241), .O(n277));
  andx  g0150(.a(n277), .b(pi14), .O(n278));
  andx  g0151(.a(n250), .b(n241), .O(n279));
  orx   g0152(.a(n279), .b(n278), .O(n280));
  andx  g0153(.a(n280), .b(n276), .O(n281));
  invx  g0154(.a(n276), .O(n282));
  andx  g0155(.a(n256), .b(n244), .O(n283));
  orx   g0156(.a(n283), .b(n243), .O(n284));
  orx   g0157(.a(n256), .b(n244), .O(n285));
  andx  g0158(.a(n285), .b(n284), .O(n286));
  andx  g0159(.a(n286), .b(n282), .O(n287));
  orx   g0160(.a(n287), .b(n281), .O(po05));
  invx  g0161(.a(pi18), .O(n289));
  andx  g0162(.a(pi19), .b(n289), .O(n290));
  invx  g0163(.a(pi19), .O(n291));
  andx  g0164(.a(n291), .b(pi18), .O(n292));
  orx   g0165(.a(n292), .b(n290), .O(n293));
  orx   g0166(.a(n267), .b(pi15), .O(n294));
  andx  g0167(.a(n294), .b(pi16), .O(n295));
  andx  g0168(.a(n267), .b(pi15), .O(n296));
  orx   g0169(.a(n296), .b(n295), .O(n297));
  andx  g0170(.a(n297), .b(n293), .O(n298));
  invx  g0171(.a(n298), .O(n299));
  orx   g0172(.a(n297), .b(n293), .O(n300));
  andx  g0173(.a(n300), .b(n299), .O(n301));
  andx  g0174(.a(n301), .b(pi20), .O(n302));
  invx  g0175(.a(pi20), .O(n303));
  invx  g0176(.a(n301), .O(n304));
  andx  g0177(.a(n304), .b(n303), .O(n305));
  orx   g0178(.a(n305), .b(n302), .O(n306));
  orx   g0179(.a(n280), .b(n271), .O(n307));
  andx  g0180(.a(n307), .b(pi17), .O(n308));
  andx  g0181(.a(n280), .b(n271), .O(n309));
  orx   g0182(.a(n309), .b(n308), .O(n310));
  andx  g0183(.a(n310), .b(n306), .O(n311));
  invx  g0184(.a(n306), .O(n312));
  andx  g0185(.a(n286), .b(n274), .O(n313));
  orx   g0186(.a(n313), .b(n273), .O(n314));
  orx   g0187(.a(n286), .b(n274), .O(n315));
  andx  g0188(.a(n315), .b(n314), .O(n316));
  andx  g0189(.a(n316), .b(n312), .O(n317));
  orx   g0190(.a(n317), .b(n311), .O(po06));
  invx  g0191(.a(pi21), .O(n319));
  andx  g0192(.a(pi22), .b(n319), .O(n320));
  invx  g0193(.a(pi22), .O(n321));
  andx  g0194(.a(n321), .b(pi21), .O(n322));
  orx   g0195(.a(n322), .b(n320), .O(n323));
  orx   g0196(.a(n297), .b(pi18), .O(n324));
  andx  g0197(.a(n324), .b(pi19), .O(n325));
  andx  g0198(.a(n297), .b(pi18), .O(n326));
  orx   g0199(.a(n326), .b(n325), .O(n327));
  andx  g0200(.a(n327), .b(n323), .O(n328));
  invx  g0201(.a(n328), .O(n329));
  orx   g0202(.a(n327), .b(n323), .O(n330));
  andx  g0203(.a(n330), .b(n329), .O(n331));
  andx  g0204(.a(n331), .b(pi23), .O(n332));
  invx  g0205(.a(pi23), .O(n333));
  invx  g0206(.a(n331), .O(n334));
  andx  g0207(.a(n334), .b(n333), .O(n335));
  orx   g0208(.a(n335), .b(n332), .O(n336));
  orx   g0209(.a(n310), .b(n301), .O(n337));
  andx  g0210(.a(n337), .b(pi20), .O(n338));
  andx  g0211(.a(n310), .b(n301), .O(n339));
  orx   g0212(.a(n339), .b(n338), .O(n340));
  andx  g0213(.a(n340), .b(n336), .O(n341));
  invx  g0214(.a(n336), .O(n342));
  andx  g0215(.a(n316), .b(n304), .O(n343));
  orx   g0216(.a(n343), .b(n303), .O(n344));
  orx   g0217(.a(n316), .b(n304), .O(n345));
  andx  g0218(.a(n345), .b(n344), .O(n346));
  andx  g0219(.a(n346), .b(n342), .O(n347));
  orx   g0220(.a(n347), .b(n341), .O(po07));
  invx  g0221(.a(pi24), .O(n349));
  andx  g0222(.a(pi25), .b(n349), .O(n350));
  invx  g0223(.a(pi25), .O(n351));
  andx  g0224(.a(n351), .b(pi24), .O(n352));
  orx   g0225(.a(n352), .b(n350), .O(n353));
  orx   g0226(.a(n327), .b(pi21), .O(n354));
  andx  g0227(.a(n354), .b(pi22), .O(n355));
  andx  g0228(.a(n327), .b(pi21), .O(n356));
  orx   g0229(.a(n356), .b(n355), .O(n357));
  andx  g0230(.a(n357), .b(n353), .O(n358));
  invx  g0231(.a(n358), .O(n359));
  orx   g0232(.a(n357), .b(n353), .O(n360));
  andx  g0233(.a(n360), .b(n359), .O(n361));
  andx  g0234(.a(n361), .b(pi26), .O(n362));
  invx  g0235(.a(pi26), .O(n363));
  invx  g0236(.a(n361), .O(n364));
  andx  g0237(.a(n364), .b(n363), .O(n365));
  orx   g0238(.a(n365), .b(n362), .O(n366));
  orx   g0239(.a(n340), .b(n331), .O(n367));
  andx  g0240(.a(n367), .b(pi23), .O(n368));
  andx  g0241(.a(n340), .b(n331), .O(n369));
  orx   g0242(.a(n369), .b(n368), .O(n370));
  andx  g0243(.a(n370), .b(n366), .O(n371));
  invx  g0244(.a(n366), .O(n372));
  andx  g0245(.a(n346), .b(n334), .O(n373));
  orx   g0246(.a(n373), .b(n333), .O(n374));
  orx   g0247(.a(n346), .b(n334), .O(n375));
  andx  g0248(.a(n375), .b(n374), .O(n376));
  andx  g0249(.a(n376), .b(n372), .O(n377));
  orx   g0250(.a(n377), .b(n371), .O(po08));
  invx  g0251(.a(pi27), .O(n379));
  andx  g0252(.a(pi28), .b(n379), .O(n380));
  invx  g0253(.a(pi28), .O(n381));
  andx  g0254(.a(n381), .b(pi27), .O(n382));
  orx   g0255(.a(n382), .b(n380), .O(n383));
  orx   g0256(.a(n357), .b(pi24), .O(n384));
  andx  g0257(.a(n384), .b(pi25), .O(n385));
  andx  g0258(.a(n357), .b(pi24), .O(n386));
  orx   g0259(.a(n386), .b(n385), .O(n387));
  andx  g0260(.a(n387), .b(n383), .O(n388));
  invx  g0261(.a(n388), .O(n389));
  orx   g0262(.a(n387), .b(n383), .O(n390));
  andx  g0263(.a(n390), .b(n389), .O(n391));
  andx  g0264(.a(n391), .b(pi29), .O(n392));
  invx  g0265(.a(pi29), .O(n393));
  invx  g0266(.a(n391), .O(n394));
  andx  g0267(.a(n394), .b(n393), .O(n395));
  orx   g0268(.a(n395), .b(n392), .O(n396));
  orx   g0269(.a(n370), .b(n361), .O(n397));
  andx  g0270(.a(n397), .b(pi26), .O(n398));
  andx  g0271(.a(n370), .b(n361), .O(n399));
  orx   g0272(.a(n399), .b(n398), .O(n400));
  andx  g0273(.a(n400), .b(n396), .O(n401));
  invx  g0274(.a(n396), .O(n402));
  andx  g0275(.a(n376), .b(n364), .O(n403));
  orx   g0276(.a(n403), .b(n363), .O(n404));
  orx   g0277(.a(n376), .b(n364), .O(n405));
  andx  g0278(.a(n405), .b(n404), .O(n406));
  andx  g0279(.a(n406), .b(n402), .O(n407));
  orx   g0280(.a(n407), .b(n401), .O(po09));
  invx  g0281(.a(pi30), .O(n409));
  andx  g0282(.a(pi31), .b(n409), .O(n410));
  invx  g0283(.a(pi31), .O(n411));
  andx  g0284(.a(n411), .b(pi30), .O(n412));
  orx   g0285(.a(n412), .b(n410), .O(n413));
  orx   g0286(.a(n387), .b(pi27), .O(n414));
  andx  g0287(.a(n414), .b(pi28), .O(n415));
  andx  g0288(.a(n387), .b(pi27), .O(n416));
  orx   g0289(.a(n416), .b(n415), .O(n417));
  andx  g0290(.a(n417), .b(n413), .O(n418));
  invx  g0291(.a(n418), .O(n419));
  orx   g0292(.a(n417), .b(n413), .O(n420));
  andx  g0293(.a(n420), .b(n419), .O(n421));
  andx  g0294(.a(n421), .b(pi32), .O(n422));
  invx  g0295(.a(pi32), .O(n423));
  invx  g0296(.a(n421), .O(n424));
  andx  g0297(.a(n424), .b(n423), .O(n425));
  orx   g0298(.a(n425), .b(n422), .O(n426));
  orx   g0299(.a(n400), .b(n391), .O(n427));
  andx  g0300(.a(n427), .b(pi29), .O(n428));
  andx  g0301(.a(n400), .b(n391), .O(n429));
  orx   g0302(.a(n429), .b(n428), .O(n430));
  andx  g0303(.a(n430), .b(n426), .O(n431));
  invx  g0304(.a(n426), .O(n432));
  andx  g0305(.a(n406), .b(n394), .O(n433));
  orx   g0306(.a(n433), .b(n393), .O(n434));
  orx   g0307(.a(n406), .b(n394), .O(n435));
  andx  g0308(.a(n435), .b(n434), .O(n436));
  andx  g0309(.a(n436), .b(n432), .O(n437));
  orx   g0310(.a(n437), .b(n431), .O(po10));
  invx  g0311(.a(pi33), .O(n439));
  andx  g0312(.a(pi34), .b(n439), .O(n440));
  invx  g0313(.a(pi34), .O(n441));
  andx  g0314(.a(n441), .b(pi33), .O(n442));
  orx   g0315(.a(n442), .b(n440), .O(n443));
  orx   g0316(.a(n417), .b(pi30), .O(n444));
  andx  g0317(.a(n444), .b(pi31), .O(n445));
  andx  g0318(.a(n417), .b(pi30), .O(n446));
  orx   g0319(.a(n446), .b(n445), .O(n447));
  andx  g0320(.a(n447), .b(n443), .O(n448));
  invx  g0321(.a(n448), .O(n449));
  orx   g0322(.a(n447), .b(n443), .O(n450));
  andx  g0323(.a(n450), .b(n449), .O(n451));
  andx  g0324(.a(n451), .b(pi35), .O(n452));
  invx  g0325(.a(pi35), .O(n453));
  invx  g0326(.a(n451), .O(n454));
  andx  g0327(.a(n454), .b(n453), .O(n455));
  orx   g0328(.a(n455), .b(n452), .O(n456));
  orx   g0329(.a(n430), .b(n421), .O(n457));
  andx  g0330(.a(n457), .b(pi32), .O(n458));
  andx  g0331(.a(n430), .b(n421), .O(n459));
  orx   g0332(.a(n459), .b(n458), .O(n460));
  andx  g0333(.a(n460), .b(n456), .O(n461));
  invx  g0334(.a(n456), .O(n462));
  andx  g0335(.a(n436), .b(n424), .O(n463));
  orx   g0336(.a(n463), .b(n423), .O(n464));
  orx   g0337(.a(n436), .b(n424), .O(n465));
  andx  g0338(.a(n465), .b(n464), .O(n466));
  andx  g0339(.a(n466), .b(n462), .O(n467));
  orx   g0340(.a(n467), .b(n461), .O(po11));
  invx  g0341(.a(pi36), .O(n469));
  andx  g0342(.a(pi37), .b(n469), .O(n470));
  invx  g0343(.a(pi37), .O(n471));
  andx  g0344(.a(n471), .b(pi36), .O(n472));
  orx   g0345(.a(n472), .b(n470), .O(n473));
  orx   g0346(.a(n447), .b(pi33), .O(n474));
  andx  g0347(.a(n474), .b(pi34), .O(n475));
  andx  g0348(.a(n447), .b(pi33), .O(n476));
  orx   g0349(.a(n476), .b(n475), .O(n477));
  andx  g0350(.a(n477), .b(n473), .O(n478));
  invx  g0351(.a(n478), .O(n479));
  orx   g0352(.a(n477), .b(n473), .O(n480));
  andx  g0353(.a(n480), .b(n479), .O(n481));
  andx  g0354(.a(n481), .b(pi38), .O(n482));
  invx  g0355(.a(pi38), .O(n483));
  invx  g0356(.a(n481), .O(n484));
  andx  g0357(.a(n484), .b(n483), .O(n485));
  orx   g0358(.a(n485), .b(n482), .O(n486));
  orx   g0359(.a(n460), .b(n451), .O(n487));
  andx  g0360(.a(n487), .b(pi35), .O(n488));
  andx  g0361(.a(n460), .b(n451), .O(n489));
  orx   g0362(.a(n489), .b(n488), .O(n490));
  andx  g0363(.a(n490), .b(n486), .O(n491));
  invx  g0364(.a(n486), .O(n492));
  andx  g0365(.a(n466), .b(n454), .O(n493));
  orx   g0366(.a(n493), .b(n453), .O(n494));
  orx   g0367(.a(n466), .b(n454), .O(n495));
  andx  g0368(.a(n495), .b(n494), .O(n496));
  andx  g0369(.a(n496), .b(n492), .O(n497));
  orx   g0370(.a(n497), .b(n491), .O(po12));
  invx  g0371(.a(pi39), .O(n499));
  andx  g0372(.a(pi40), .b(n499), .O(n500));
  invx  g0373(.a(pi40), .O(n501));
  andx  g0374(.a(n501), .b(pi39), .O(n502));
  orx   g0375(.a(n502), .b(n500), .O(n503));
  orx   g0376(.a(n477), .b(pi36), .O(n504));
  andx  g0377(.a(n504), .b(pi37), .O(n505));
  andx  g0378(.a(n477), .b(pi36), .O(n506));
  orx   g0379(.a(n506), .b(n505), .O(n507));
  andx  g0380(.a(n507), .b(n503), .O(n508));
  invx  g0381(.a(n508), .O(n509));
  orx   g0382(.a(n507), .b(n503), .O(n510));
  andx  g0383(.a(n510), .b(n509), .O(n511));
  andx  g0384(.a(n511), .b(pi41), .O(n512));
  invx  g0385(.a(pi41), .O(n513));
  invx  g0386(.a(n511), .O(n514));
  andx  g0387(.a(n514), .b(n513), .O(n515));
  orx   g0388(.a(n515), .b(n512), .O(n516));
  orx   g0389(.a(n490), .b(n481), .O(n517));
  andx  g0390(.a(n517), .b(pi38), .O(n518));
  andx  g0391(.a(n490), .b(n481), .O(n519));
  orx   g0392(.a(n519), .b(n518), .O(n520));
  andx  g0393(.a(n520), .b(n516), .O(n521));
  invx  g0394(.a(n516), .O(n522));
  andx  g0395(.a(n496), .b(n484), .O(n523));
  orx   g0396(.a(n523), .b(n483), .O(n524));
  orx   g0397(.a(n496), .b(n484), .O(n525));
  andx  g0398(.a(n525), .b(n524), .O(n526));
  andx  g0399(.a(n526), .b(n522), .O(n527));
  orx   g0400(.a(n527), .b(n521), .O(po13));
  invx  g0401(.a(pi42), .O(n529));
  andx  g0402(.a(pi43), .b(n529), .O(n530));
  invx  g0403(.a(pi43), .O(n531));
  andx  g0404(.a(n531), .b(pi42), .O(n532));
  orx   g0405(.a(n532), .b(n530), .O(n533));
  orx   g0406(.a(n507), .b(pi39), .O(n534));
  andx  g0407(.a(n534), .b(pi40), .O(n535));
  andx  g0408(.a(n507), .b(pi39), .O(n536));
  orx   g0409(.a(n536), .b(n535), .O(n537));
  andx  g0410(.a(n537), .b(n533), .O(n538));
  invx  g0411(.a(n538), .O(n539));
  orx   g0412(.a(n537), .b(n533), .O(n540));
  andx  g0413(.a(n540), .b(n539), .O(n541));
  andx  g0414(.a(n541), .b(pi44), .O(n542));
  invx  g0415(.a(pi44), .O(n543));
  invx  g0416(.a(n541), .O(n544));
  andx  g0417(.a(n544), .b(n543), .O(n545));
  orx   g0418(.a(n545), .b(n542), .O(n546));
  orx   g0419(.a(n520), .b(n511), .O(n547));
  andx  g0420(.a(n547), .b(pi41), .O(n548));
  andx  g0421(.a(n520), .b(n511), .O(n549));
  orx   g0422(.a(n549), .b(n548), .O(n550));
  andx  g0423(.a(n550), .b(n546), .O(n551));
  invx  g0424(.a(n546), .O(n552));
  andx  g0425(.a(n526), .b(n514), .O(n553));
  orx   g0426(.a(n553), .b(n513), .O(n554));
  orx   g0427(.a(n526), .b(n514), .O(n555));
  andx  g0428(.a(n555), .b(n554), .O(n556));
  andx  g0429(.a(n556), .b(n552), .O(n557));
  orx   g0430(.a(n557), .b(n551), .O(po14));
  invx  g0431(.a(pi45), .O(n559));
  andx  g0432(.a(pi46), .b(n559), .O(n560));
  invx  g0433(.a(pi46), .O(n561));
  andx  g0434(.a(n561), .b(pi45), .O(n562));
  orx   g0435(.a(n562), .b(n560), .O(n563));
  orx   g0436(.a(n537), .b(pi42), .O(n564));
  andx  g0437(.a(n564), .b(pi43), .O(n565));
  andx  g0438(.a(n537), .b(pi42), .O(n566));
  orx   g0439(.a(n566), .b(n565), .O(n567));
  andx  g0440(.a(n567), .b(n563), .O(n568));
  invx  g0441(.a(n568), .O(n569));
  orx   g0442(.a(n567), .b(n563), .O(n570));
  andx  g0443(.a(n570), .b(n569), .O(n571));
  andx  g0444(.a(n571), .b(pi47), .O(n572));
  invx  g0445(.a(pi47), .O(n573));
  invx  g0446(.a(n571), .O(n574));
  andx  g0447(.a(n574), .b(n573), .O(n575));
  orx   g0448(.a(n575), .b(n572), .O(n576));
  orx   g0449(.a(n550), .b(n541), .O(n577));
  andx  g0450(.a(n577), .b(pi44), .O(n578));
  andx  g0451(.a(n550), .b(n541), .O(n579));
  orx   g0452(.a(n579), .b(n578), .O(n580));
  andx  g0453(.a(n580), .b(n576), .O(n581));
  invx  g0454(.a(n576), .O(n582));
  andx  g0455(.a(n556), .b(n544), .O(n583));
  orx   g0456(.a(n583), .b(n543), .O(n584));
  orx   g0457(.a(n556), .b(n544), .O(n585));
  andx  g0458(.a(n585), .b(n584), .O(n586));
  andx  g0459(.a(n586), .b(n582), .O(n587));
  orx   g0460(.a(n587), .b(n581), .O(po15));
  invx  g0461(.a(pi48), .O(n589));
  andx  g0462(.a(pi49), .b(n589), .O(n590));
  invx  g0463(.a(pi49), .O(n591));
  andx  g0464(.a(n591), .b(pi48), .O(n592));
  orx   g0465(.a(n592), .b(n590), .O(n593));
  orx   g0466(.a(n567), .b(pi45), .O(n594));
  andx  g0467(.a(n594), .b(pi46), .O(n595));
  andx  g0468(.a(n567), .b(pi45), .O(n596));
  orx   g0469(.a(n596), .b(n595), .O(n597));
  andx  g0470(.a(n597), .b(n593), .O(n598));
  invx  g0471(.a(n598), .O(n599));
  orx   g0472(.a(n597), .b(n593), .O(n600));
  andx  g0473(.a(n600), .b(n599), .O(n601));
  andx  g0474(.a(n601), .b(pi50), .O(n602));
  invx  g0475(.a(pi50), .O(n603));
  invx  g0476(.a(n601), .O(n604));
  andx  g0477(.a(n604), .b(n603), .O(n605));
  orx   g0478(.a(n605), .b(n602), .O(n606));
  orx   g0479(.a(n580), .b(n571), .O(n607));
  andx  g0480(.a(n607), .b(pi47), .O(n608));
  andx  g0481(.a(n580), .b(n571), .O(n609));
  orx   g0482(.a(n609), .b(n608), .O(n610));
  andx  g0483(.a(n610), .b(n606), .O(n611));
  invx  g0484(.a(n606), .O(n612));
  andx  g0485(.a(n586), .b(n574), .O(n613));
  orx   g0486(.a(n613), .b(n573), .O(n614));
  orx   g0487(.a(n586), .b(n574), .O(n615));
  andx  g0488(.a(n615), .b(n614), .O(n616));
  andx  g0489(.a(n616), .b(n612), .O(n617));
  orx   g0490(.a(n617), .b(n611), .O(po16));
  invx  g0491(.a(pi51), .O(n619));
  andx  g0492(.a(pi52), .b(n619), .O(n620));
  invx  g0493(.a(pi52), .O(n621));
  andx  g0494(.a(n621), .b(pi51), .O(n622));
  orx   g0495(.a(n622), .b(n620), .O(n623));
  orx   g0496(.a(n597), .b(pi48), .O(n624));
  andx  g0497(.a(n624), .b(pi49), .O(n625));
  andx  g0498(.a(n597), .b(pi48), .O(n626));
  orx   g0499(.a(n626), .b(n625), .O(n627));
  andx  g0500(.a(n627), .b(n623), .O(n628));
  invx  g0501(.a(n628), .O(n629));
  orx   g0502(.a(n627), .b(n623), .O(n630));
  andx  g0503(.a(n630), .b(n629), .O(n631));
  andx  g0504(.a(n631), .b(pi53), .O(n632));
  invx  g0505(.a(pi53), .O(n633));
  invx  g0506(.a(n631), .O(n634));
  andx  g0507(.a(n634), .b(n633), .O(n635));
  orx   g0508(.a(n635), .b(n632), .O(n636));
  orx   g0509(.a(n610), .b(n601), .O(n637));
  andx  g0510(.a(n637), .b(pi50), .O(n638));
  andx  g0511(.a(n610), .b(n601), .O(n639));
  orx   g0512(.a(n639), .b(n638), .O(n640));
  andx  g0513(.a(n640), .b(n636), .O(n641));
  invx  g0514(.a(n636), .O(n642));
  andx  g0515(.a(n616), .b(n604), .O(n643));
  orx   g0516(.a(n643), .b(n603), .O(n644));
  orx   g0517(.a(n616), .b(n604), .O(n645));
  andx  g0518(.a(n645), .b(n644), .O(n646));
  andx  g0519(.a(n646), .b(n642), .O(n647));
  orx   g0520(.a(n647), .b(n641), .O(po17));
  invx  g0521(.a(pi54), .O(n649));
  andx  g0522(.a(pi55), .b(n649), .O(n650));
  invx  g0523(.a(pi55), .O(n651));
  andx  g0524(.a(n651), .b(pi54), .O(n652));
  orx   g0525(.a(n652), .b(n650), .O(n653));
  orx   g0526(.a(n627), .b(pi51), .O(n654));
  andx  g0527(.a(n654), .b(pi52), .O(n655));
  andx  g0528(.a(n627), .b(pi51), .O(n656));
  orx   g0529(.a(n656), .b(n655), .O(n657));
  andx  g0530(.a(n657), .b(n653), .O(n658));
  invx  g0531(.a(n658), .O(n659));
  orx   g0532(.a(n657), .b(n653), .O(n660));
  andx  g0533(.a(n660), .b(n659), .O(n661));
  andx  g0534(.a(n661), .b(pi56), .O(n662));
  invx  g0535(.a(pi56), .O(n663));
  invx  g0536(.a(n661), .O(n664));
  andx  g0537(.a(n664), .b(n663), .O(n665));
  orx   g0538(.a(n665), .b(n662), .O(n666));
  orx   g0539(.a(n640), .b(n631), .O(n667));
  andx  g0540(.a(n667), .b(pi53), .O(n668));
  andx  g0541(.a(n640), .b(n631), .O(n669));
  orx   g0542(.a(n669), .b(n668), .O(n670));
  andx  g0543(.a(n670), .b(n666), .O(n671));
  invx  g0544(.a(n666), .O(n672));
  andx  g0545(.a(n646), .b(n634), .O(n673));
  orx   g0546(.a(n673), .b(n633), .O(n674));
  orx   g0547(.a(n646), .b(n634), .O(n675));
  andx  g0548(.a(n675), .b(n674), .O(n676));
  andx  g0549(.a(n676), .b(n672), .O(n677));
  orx   g0550(.a(n677), .b(n671), .O(po18));
  invx  g0551(.a(pi57), .O(n679));
  andx  g0552(.a(pi58), .b(n679), .O(n680));
  invx  g0553(.a(pi58), .O(n681));
  andx  g0554(.a(n681), .b(pi57), .O(n682));
  orx   g0555(.a(n682), .b(n680), .O(n683));
  orx   g0556(.a(n657), .b(pi54), .O(n684));
  andx  g0557(.a(n684), .b(pi55), .O(n685));
  andx  g0558(.a(n657), .b(pi54), .O(n686));
  orx   g0559(.a(n686), .b(n685), .O(n687));
  andx  g0560(.a(n687), .b(n683), .O(n688));
  invx  g0561(.a(n688), .O(n689));
  orx   g0562(.a(n687), .b(n683), .O(n690));
  andx  g0563(.a(n690), .b(n689), .O(n691));
  andx  g0564(.a(n691), .b(pi59), .O(n692));
  invx  g0565(.a(pi59), .O(n693));
  invx  g0566(.a(n691), .O(n694));
  andx  g0567(.a(n694), .b(n693), .O(n695));
  orx   g0568(.a(n695), .b(n692), .O(n696));
  orx   g0569(.a(n670), .b(n661), .O(n697));
  andx  g0570(.a(n697), .b(pi56), .O(n698));
  andx  g0571(.a(n670), .b(n661), .O(n699));
  orx   g0572(.a(n699), .b(n698), .O(n700));
  andx  g0573(.a(n700), .b(n696), .O(n701));
  invx  g0574(.a(n696), .O(n702));
  andx  g0575(.a(n676), .b(n664), .O(n703));
  orx   g0576(.a(n703), .b(n663), .O(n704));
  orx   g0577(.a(n676), .b(n664), .O(n705));
  andx  g0578(.a(n705), .b(n704), .O(n706));
  andx  g0579(.a(n706), .b(n702), .O(n707));
  orx   g0580(.a(n707), .b(n701), .O(po19));
  invx  g0581(.a(pi60), .O(n709));
  andx  g0582(.a(pi61), .b(n709), .O(n710));
  invx  g0583(.a(pi61), .O(n711));
  andx  g0584(.a(n711), .b(pi60), .O(n712));
  orx   g0585(.a(n712), .b(n710), .O(n713));
  orx   g0586(.a(n687), .b(pi57), .O(n714));
  andx  g0587(.a(n714), .b(pi58), .O(n715));
  andx  g0588(.a(n687), .b(pi57), .O(n716));
  orx   g0589(.a(n716), .b(n715), .O(n717));
  andx  g0590(.a(n717), .b(n713), .O(n718));
  invx  g0591(.a(n718), .O(n719));
  orx   g0592(.a(n717), .b(n713), .O(n720));
  andx  g0593(.a(n720), .b(n719), .O(n721));
  andx  g0594(.a(n721), .b(pi62), .O(n722));
  invx  g0595(.a(pi62), .O(n723));
  invx  g0596(.a(n721), .O(n724));
  andx  g0597(.a(n724), .b(n723), .O(n725));
  orx   g0598(.a(n725), .b(n722), .O(n726));
  orx   g0599(.a(n700), .b(n691), .O(n727));
  andx  g0600(.a(n727), .b(pi59), .O(n728));
  andx  g0601(.a(n700), .b(n691), .O(n729));
  orx   g0602(.a(n729), .b(n728), .O(n730));
  andx  g0603(.a(n730), .b(n726), .O(n731));
  invx  g0604(.a(n726), .O(n732));
  andx  g0605(.a(n706), .b(n694), .O(n733));
  orx   g0606(.a(n733), .b(n693), .O(n734));
  orx   g0607(.a(n706), .b(n694), .O(n735));
  andx  g0608(.a(n735), .b(n734), .O(n736));
  andx  g0609(.a(n736), .b(n732), .O(n737));
  orx   g0610(.a(n737), .b(n731), .O(po20));
  invx  g0611(.a(pi63), .O(n739));
  andx  g0612(.a(pi64), .b(n739), .O(n740));
  invx  g0613(.a(pi64), .O(n741));
  andx  g0614(.a(n741), .b(pi63), .O(n742));
  orx   g0615(.a(n742), .b(n740), .O(n743));
  orx   g0616(.a(n717), .b(pi60), .O(n744));
  andx  g0617(.a(n744), .b(pi61), .O(n745));
  andx  g0618(.a(n717), .b(pi60), .O(n746));
  orx   g0619(.a(n746), .b(n745), .O(n747));
  andx  g0620(.a(n747), .b(n743), .O(n748));
  invx  g0621(.a(n748), .O(n749));
  orx   g0622(.a(n747), .b(n743), .O(n750));
  andx  g0623(.a(n750), .b(n749), .O(n751));
  andx  g0624(.a(n751), .b(pi65), .O(n752));
  invx  g0625(.a(pi65), .O(n753));
  invx  g0626(.a(n751), .O(n754));
  andx  g0627(.a(n754), .b(n753), .O(n755));
  orx   g0628(.a(n755), .b(n752), .O(n756));
  orx   g0629(.a(n730), .b(n721), .O(n757));
  andx  g0630(.a(n757), .b(pi62), .O(n758));
  andx  g0631(.a(n730), .b(n721), .O(n759));
  orx   g0632(.a(n759), .b(n758), .O(n760));
  andx  g0633(.a(n760), .b(n756), .O(n761));
  invx  g0634(.a(n756), .O(n762));
  andx  g0635(.a(n736), .b(n724), .O(n763));
  orx   g0636(.a(n763), .b(n723), .O(n764));
  orx   g0637(.a(n736), .b(n724), .O(n765));
  andx  g0638(.a(n765), .b(n764), .O(n766));
  andx  g0639(.a(n766), .b(n762), .O(n767));
  orx   g0640(.a(n767), .b(n761), .O(po21));
  invx  g0641(.a(pi66), .O(n769));
  andx  g0642(.a(pi67), .b(n769), .O(n770));
  invx  g0643(.a(pi67), .O(n771));
  andx  g0644(.a(n771), .b(pi66), .O(n772));
  orx   g0645(.a(n772), .b(n770), .O(n773));
  orx   g0646(.a(n747), .b(pi63), .O(n774));
  andx  g0647(.a(n774), .b(pi64), .O(n775));
  andx  g0648(.a(n747), .b(pi63), .O(n776));
  orx   g0649(.a(n776), .b(n775), .O(n777));
  andx  g0650(.a(n777), .b(n773), .O(n778));
  invx  g0651(.a(n778), .O(n779));
  orx   g0652(.a(n777), .b(n773), .O(n780));
  andx  g0653(.a(n780), .b(n779), .O(n781));
  andx  g0654(.a(n781), .b(pi68), .O(n782));
  invx  g0655(.a(pi68), .O(n783));
  invx  g0656(.a(n781), .O(n784));
  andx  g0657(.a(n784), .b(n783), .O(n785));
  orx   g0658(.a(n785), .b(n782), .O(n786));
  orx   g0659(.a(n760), .b(n751), .O(n787));
  andx  g0660(.a(n787), .b(pi65), .O(n788));
  andx  g0661(.a(n760), .b(n751), .O(n789));
  orx   g0662(.a(n789), .b(n788), .O(n790));
  andx  g0663(.a(n790), .b(n786), .O(n791));
  invx  g0664(.a(n786), .O(n792));
  andx  g0665(.a(n766), .b(n754), .O(n793));
  orx   g0666(.a(n793), .b(n753), .O(n794));
  orx   g0667(.a(n766), .b(n754), .O(n795));
  andx  g0668(.a(n795), .b(n794), .O(n796));
  andx  g0669(.a(n796), .b(n792), .O(n797));
  orx   g0670(.a(n797), .b(n791), .O(po22));
  invx  g0671(.a(pi69), .O(n799));
  andx  g0672(.a(pi70), .b(n799), .O(n800));
  invx  g0673(.a(pi70), .O(n801));
  andx  g0674(.a(n801), .b(pi69), .O(n802));
  orx   g0675(.a(n802), .b(n800), .O(n803));
  orx   g0676(.a(n777), .b(pi66), .O(n804));
  andx  g0677(.a(n804), .b(pi67), .O(n805));
  andx  g0678(.a(n777), .b(pi66), .O(n806));
  orx   g0679(.a(n806), .b(n805), .O(n807));
  andx  g0680(.a(n807), .b(n803), .O(n808));
  invx  g0681(.a(n808), .O(n809));
  orx   g0682(.a(n807), .b(n803), .O(n810));
  andx  g0683(.a(n810), .b(n809), .O(n811));
  andx  g0684(.a(n811), .b(pi71), .O(n812));
  invx  g0685(.a(pi71), .O(n813));
  invx  g0686(.a(n811), .O(n814));
  andx  g0687(.a(n814), .b(n813), .O(n815));
  orx   g0688(.a(n815), .b(n812), .O(n816));
  orx   g0689(.a(n790), .b(n781), .O(n817));
  andx  g0690(.a(n817), .b(pi68), .O(n818));
  andx  g0691(.a(n790), .b(n781), .O(n819));
  orx   g0692(.a(n819), .b(n818), .O(n820));
  andx  g0693(.a(n820), .b(n816), .O(n821));
  invx  g0694(.a(n816), .O(n822));
  andx  g0695(.a(n796), .b(n784), .O(n823));
  orx   g0696(.a(n823), .b(n783), .O(n824));
  orx   g0697(.a(n796), .b(n784), .O(n825));
  andx  g0698(.a(n825), .b(n824), .O(n826));
  andx  g0699(.a(n826), .b(n822), .O(n827));
  orx   g0700(.a(n827), .b(n821), .O(po23));
  invx  g0701(.a(pi72), .O(n829));
  andx  g0702(.a(pi73), .b(n829), .O(n830));
  invx  g0703(.a(pi73), .O(n831));
  andx  g0704(.a(n831), .b(pi72), .O(n832));
  orx   g0705(.a(n832), .b(n830), .O(n833));
  orx   g0706(.a(n807), .b(pi69), .O(n834));
  andx  g0707(.a(n834), .b(pi70), .O(n835));
  andx  g0708(.a(n807), .b(pi69), .O(n836));
  orx   g0709(.a(n836), .b(n835), .O(n837));
  andx  g0710(.a(n837), .b(n833), .O(n838));
  invx  g0711(.a(n838), .O(n839));
  orx   g0712(.a(n837), .b(n833), .O(n840));
  andx  g0713(.a(n840), .b(n839), .O(n841));
  andx  g0714(.a(n841), .b(pi74), .O(n842));
  invx  g0715(.a(pi74), .O(n843));
  invx  g0716(.a(n841), .O(n844));
  andx  g0717(.a(n844), .b(n843), .O(n845));
  orx   g0718(.a(n845), .b(n842), .O(n846));
  orx   g0719(.a(n820), .b(n811), .O(n847));
  andx  g0720(.a(n847), .b(pi71), .O(n848));
  andx  g0721(.a(n820), .b(n811), .O(n849));
  orx   g0722(.a(n849), .b(n848), .O(n850));
  andx  g0723(.a(n850), .b(n846), .O(n851));
  invx  g0724(.a(n846), .O(n852));
  andx  g0725(.a(n826), .b(n814), .O(n853));
  orx   g0726(.a(n853), .b(n813), .O(n854));
  orx   g0727(.a(n826), .b(n814), .O(n855));
  andx  g0728(.a(n855), .b(n854), .O(n856));
  andx  g0729(.a(n856), .b(n852), .O(n857));
  orx   g0730(.a(n857), .b(n851), .O(po24));
  invx  g0731(.a(pi75), .O(n859));
  andx  g0732(.a(pi76), .b(n859), .O(n860));
  invx  g0733(.a(pi76), .O(n861));
  andx  g0734(.a(n861), .b(pi75), .O(n862));
  orx   g0735(.a(n862), .b(n860), .O(n863));
  orx   g0736(.a(n837), .b(pi72), .O(n864));
  andx  g0737(.a(n864), .b(pi73), .O(n865));
  andx  g0738(.a(n837), .b(pi72), .O(n866));
  orx   g0739(.a(n866), .b(n865), .O(n867));
  andx  g0740(.a(n867), .b(n863), .O(n868));
  invx  g0741(.a(n868), .O(n869));
  orx   g0742(.a(n867), .b(n863), .O(n870));
  andx  g0743(.a(n870), .b(n869), .O(n871));
  andx  g0744(.a(n871), .b(pi77), .O(n872));
  invx  g0745(.a(pi77), .O(n873));
  invx  g0746(.a(n871), .O(n874));
  andx  g0747(.a(n874), .b(n873), .O(n875));
  orx   g0748(.a(n875), .b(n872), .O(n876));
  orx   g0749(.a(n850), .b(n841), .O(n877));
  andx  g0750(.a(n877), .b(pi74), .O(n878));
  andx  g0751(.a(n850), .b(n841), .O(n879));
  orx   g0752(.a(n879), .b(n878), .O(n880));
  andx  g0753(.a(n880), .b(n876), .O(n881));
  invx  g0754(.a(n876), .O(n882));
  andx  g0755(.a(n856), .b(n844), .O(n883));
  orx   g0756(.a(n883), .b(n843), .O(n884));
  orx   g0757(.a(n856), .b(n844), .O(n885));
  andx  g0758(.a(n885), .b(n884), .O(n886));
  andx  g0759(.a(n886), .b(n882), .O(n887));
  orx   g0760(.a(n887), .b(n881), .O(po25));
  invx  g0761(.a(pi78), .O(n889));
  andx  g0762(.a(pi79), .b(n889), .O(n890));
  invx  g0763(.a(pi79), .O(n891));
  andx  g0764(.a(n891), .b(pi78), .O(n892));
  orx   g0765(.a(n892), .b(n890), .O(n893));
  orx   g0766(.a(n867), .b(pi75), .O(n894));
  andx  g0767(.a(n894), .b(pi76), .O(n895));
  andx  g0768(.a(n867), .b(pi75), .O(n896));
  orx   g0769(.a(n896), .b(n895), .O(n897));
  andx  g0770(.a(n897), .b(n893), .O(n898));
  invx  g0771(.a(n898), .O(n899));
  orx   g0772(.a(n897), .b(n893), .O(n900));
  andx  g0773(.a(n900), .b(n899), .O(n901));
  andx  g0774(.a(n901), .b(pi80), .O(n902));
  invx  g0775(.a(pi80), .O(n903));
  invx  g0776(.a(n901), .O(n904));
  andx  g0777(.a(n904), .b(n903), .O(n905));
  orx   g0778(.a(n905), .b(n902), .O(n906));
  orx   g0779(.a(n880), .b(n871), .O(n907));
  andx  g0780(.a(n907), .b(pi77), .O(n908));
  andx  g0781(.a(n880), .b(n871), .O(n909));
  orx   g0782(.a(n909), .b(n908), .O(n910));
  andx  g0783(.a(n910), .b(n906), .O(n911));
  invx  g0784(.a(n906), .O(n912));
  andx  g0785(.a(n886), .b(n874), .O(n913));
  orx   g0786(.a(n913), .b(n873), .O(n914));
  orx   g0787(.a(n886), .b(n874), .O(n915));
  andx  g0788(.a(n915), .b(n914), .O(n916));
  andx  g0789(.a(n916), .b(n912), .O(n917));
  orx   g0790(.a(n917), .b(n911), .O(po26));
  invx  g0791(.a(pi81), .O(n919));
  andx  g0792(.a(pi82), .b(n919), .O(n920));
  invx  g0793(.a(pi82), .O(n921));
  andx  g0794(.a(n921), .b(pi81), .O(n922));
  orx   g0795(.a(n922), .b(n920), .O(n923));
  orx   g0796(.a(n897), .b(pi78), .O(n924));
  andx  g0797(.a(n924), .b(pi79), .O(n925));
  andx  g0798(.a(n897), .b(pi78), .O(n926));
  orx   g0799(.a(n926), .b(n925), .O(n927));
  andx  g0800(.a(n927), .b(n923), .O(n928));
  invx  g0801(.a(n928), .O(n929));
  orx   g0802(.a(n927), .b(n923), .O(n930));
  andx  g0803(.a(n930), .b(n929), .O(n931));
  andx  g0804(.a(n931), .b(pi83), .O(n932));
  invx  g0805(.a(pi83), .O(n933));
  invx  g0806(.a(n931), .O(n934));
  andx  g0807(.a(n934), .b(n933), .O(n935));
  orx   g0808(.a(n935), .b(n932), .O(n936));
  orx   g0809(.a(n910), .b(n901), .O(n937));
  andx  g0810(.a(n937), .b(pi80), .O(n938));
  andx  g0811(.a(n910), .b(n901), .O(n939));
  orx   g0812(.a(n939), .b(n938), .O(n940));
  andx  g0813(.a(n940), .b(n936), .O(n941));
  invx  g0814(.a(n936), .O(n942));
  andx  g0815(.a(n916), .b(n904), .O(n943));
  orx   g0816(.a(n943), .b(n903), .O(n944));
  orx   g0817(.a(n916), .b(n904), .O(n945));
  andx  g0818(.a(n945), .b(n944), .O(n946));
  andx  g0819(.a(n946), .b(n942), .O(n947));
  orx   g0820(.a(n947), .b(n941), .O(po27));
  invx  g0821(.a(pi84), .O(n949));
  andx  g0822(.a(pi85), .b(n949), .O(n950));
  invx  g0823(.a(pi85), .O(n951));
  andx  g0824(.a(n951), .b(pi84), .O(n952));
  orx   g0825(.a(n952), .b(n950), .O(n953));
  orx   g0826(.a(n927), .b(pi81), .O(n954));
  andx  g0827(.a(n954), .b(pi82), .O(n955));
  andx  g0828(.a(n927), .b(pi81), .O(n956));
  orx   g0829(.a(n956), .b(n955), .O(n957));
  andx  g0830(.a(n957), .b(n953), .O(n958));
  invx  g0831(.a(n958), .O(n959));
  orx   g0832(.a(n957), .b(n953), .O(n960));
  andx  g0833(.a(n960), .b(n959), .O(n961));
  andx  g0834(.a(n961), .b(pi86), .O(n962));
  invx  g0835(.a(pi86), .O(n963));
  invx  g0836(.a(n961), .O(n964));
  andx  g0837(.a(n964), .b(n963), .O(n965));
  orx   g0838(.a(n965), .b(n962), .O(n966));
  orx   g0839(.a(n940), .b(n931), .O(n967));
  andx  g0840(.a(n967), .b(pi83), .O(n968));
  andx  g0841(.a(n940), .b(n931), .O(n969));
  orx   g0842(.a(n969), .b(n968), .O(n970));
  andx  g0843(.a(n970), .b(n966), .O(n971));
  invx  g0844(.a(n966), .O(n972));
  andx  g0845(.a(n946), .b(n934), .O(n973));
  orx   g0846(.a(n973), .b(n933), .O(n974));
  orx   g0847(.a(n946), .b(n934), .O(n975));
  andx  g0848(.a(n975), .b(n974), .O(n976));
  andx  g0849(.a(n976), .b(n972), .O(n977));
  orx   g0850(.a(n977), .b(n971), .O(po28));
  invx  g0851(.a(pi87), .O(n979));
  andx  g0852(.a(pi88), .b(n979), .O(n980));
  invx  g0853(.a(pi88), .O(n981));
  andx  g0854(.a(n981), .b(pi87), .O(n982));
  orx   g0855(.a(n982), .b(n980), .O(n983));
  orx   g0856(.a(n957), .b(pi84), .O(n984));
  andx  g0857(.a(n984), .b(pi85), .O(n985));
  andx  g0858(.a(n957), .b(pi84), .O(n986));
  orx   g0859(.a(n986), .b(n985), .O(n987));
  andx  g0860(.a(n987), .b(n983), .O(n988));
  invx  g0861(.a(n988), .O(n989));
  orx   g0862(.a(n987), .b(n983), .O(n990));
  andx  g0863(.a(n990), .b(n989), .O(n991));
  andx  g0864(.a(n991), .b(pi89), .O(n992));
  invx  g0865(.a(pi89), .O(n993));
  invx  g0866(.a(n991), .O(n994));
  andx  g0867(.a(n994), .b(n993), .O(n995));
  orx   g0868(.a(n995), .b(n992), .O(n996));
  orx   g0869(.a(n970), .b(n961), .O(n997));
  andx  g0870(.a(n997), .b(pi86), .O(n998));
  andx  g0871(.a(n970), .b(n961), .O(n999));
  orx   g0872(.a(n999), .b(n998), .O(n1000));
  andx  g0873(.a(n1000), .b(n996), .O(n1001));
  invx  g0874(.a(n996), .O(n1002));
  andx  g0875(.a(n976), .b(n964), .O(n1003));
  orx   g0876(.a(n1003), .b(n963), .O(n1004));
  orx   g0877(.a(n976), .b(n964), .O(n1005));
  andx  g0878(.a(n1005), .b(n1004), .O(n1006));
  andx  g0879(.a(n1006), .b(n1002), .O(n1007));
  orx   g0880(.a(n1007), .b(n1001), .O(po29));
  invx  g0881(.a(pi90), .O(n1009));
  andx  g0882(.a(pi91), .b(n1009), .O(n1010));
  invx  g0883(.a(pi91), .O(n1011));
  andx  g0884(.a(n1011), .b(pi90), .O(n1012));
  orx   g0885(.a(n1012), .b(n1010), .O(n1013));
  orx   g0886(.a(n987), .b(pi87), .O(n1014));
  andx  g0887(.a(n1014), .b(pi88), .O(n1015));
  andx  g0888(.a(n987), .b(pi87), .O(n1016));
  orx   g0889(.a(n1016), .b(n1015), .O(n1017));
  andx  g0890(.a(n1017), .b(n1013), .O(n1018));
  invx  g0891(.a(n1018), .O(n1019));
  orx   g0892(.a(n1017), .b(n1013), .O(n1020));
  andx  g0893(.a(n1020), .b(n1019), .O(n1021));
  andx  g0894(.a(n1021), .b(pi92), .O(n1022));
  invx  g0895(.a(pi92), .O(n1023));
  invx  g0896(.a(n1021), .O(n1024));
  andx  g0897(.a(n1024), .b(n1023), .O(n1025));
  orx   g0898(.a(n1025), .b(n1022), .O(n1026));
  orx   g0899(.a(n1000), .b(n991), .O(n1027));
  andx  g0900(.a(n1027), .b(pi89), .O(n1028));
  andx  g0901(.a(n1000), .b(n991), .O(n1029));
  orx   g0902(.a(n1029), .b(n1028), .O(n1030));
  andx  g0903(.a(n1030), .b(n1026), .O(n1031));
  invx  g0904(.a(n1026), .O(n1032));
  andx  g0905(.a(n1006), .b(n994), .O(n1033));
  orx   g0906(.a(n1033), .b(n993), .O(n1034));
  orx   g0907(.a(n1006), .b(n994), .O(n1035));
  andx  g0908(.a(n1035), .b(n1034), .O(n1036));
  andx  g0909(.a(n1036), .b(n1032), .O(n1037));
  orx   g0910(.a(n1037), .b(n1031), .O(po30));
  invx  g0911(.a(pi93), .O(n1039));
  andx  g0912(.a(pi94), .b(n1039), .O(n1040));
  invx  g0913(.a(n1040), .O(n1041));
  orx   g0914(.a(pi94), .b(n1039), .O(n1042));
  andx  g0915(.a(n1042), .b(n1041), .O(n1043));
  invx  g0916(.a(n1043), .O(n1044));
  orx   g0917(.a(n1017), .b(pi90), .O(n1045));
  andx  g0918(.a(n1045), .b(pi91), .O(n1046));
  andx  g0919(.a(n1017), .b(pi90), .O(n1047));
  orx   g0920(.a(n1047), .b(n1046), .O(n1048));
  orx   g0921(.a(n1048), .b(n1044), .O(n1049));
  andx  g0922(.a(n139), .b(n138), .O(n1050));
  orx   g0923(.a(n1050), .b(n141), .O(n1051));
  andx  g0924(.a(n1051), .b(n160), .O(n1052));
  andx  g0925(.a(n1052), .b(n172), .O(n1053));
  orx   g0926(.a(n1053), .b(n174), .O(n1054));
  invx  g0927(.a(n206), .O(n1055));
  andx  g0928(.a(n1055), .b(n1054), .O(n1056));
  andx  g0929(.a(n1056), .b(n199), .O(n1057));
  orx   g0930(.a(n1057), .b(n201), .O(n1058));
  invx  g0931(.a(n236), .O(n1059));
  andx  g0932(.a(n1059), .b(n1058), .O(n1060));
  andx  g0933(.a(n1060), .b(n229), .O(n1061));
  orx   g0934(.a(n1061), .b(n231), .O(n1062));
  invx  g0935(.a(n266), .O(n1063));
  andx  g0936(.a(n1063), .b(n1062), .O(n1064));
  andx  g0937(.a(n1064), .b(n259), .O(n1065));
  orx   g0938(.a(n1065), .b(n261), .O(n1066));
  invx  g0939(.a(n296), .O(n1067));
  andx  g0940(.a(n1067), .b(n1066), .O(n1068));
  andx  g0941(.a(n1068), .b(n289), .O(n1069));
  orx   g0942(.a(n1069), .b(n291), .O(n1070));
  invx  g0943(.a(n326), .O(n1071));
  andx  g0944(.a(n1071), .b(n1070), .O(n1072));
  andx  g0945(.a(n1072), .b(n319), .O(n1073));
  orx   g0946(.a(n1073), .b(n321), .O(n1074));
  invx  g0947(.a(n356), .O(n1075));
  andx  g0948(.a(n1075), .b(n1074), .O(n1076));
  andx  g0949(.a(n1076), .b(n349), .O(n1077));
  orx   g0950(.a(n1077), .b(n351), .O(n1078));
  invx  g0951(.a(n386), .O(n1079));
  andx  g0952(.a(n1079), .b(n1078), .O(n1080));
  andx  g0953(.a(n1080), .b(n379), .O(n1081));
  orx   g0954(.a(n1081), .b(n381), .O(n1082));
  invx  g0955(.a(n416), .O(n1083));
  andx  g0956(.a(n1083), .b(n1082), .O(n1084));
  andx  g0957(.a(n1084), .b(n409), .O(n1085));
  orx   g0958(.a(n1085), .b(n411), .O(n1086));
  invx  g0959(.a(n446), .O(n1087));
  andx  g0960(.a(n1087), .b(n1086), .O(n1088));
  andx  g0961(.a(n1088), .b(n439), .O(n1089));
  orx   g0962(.a(n1089), .b(n441), .O(n1090));
  invx  g0963(.a(n476), .O(n1091));
  andx  g0964(.a(n1091), .b(n1090), .O(n1092));
  andx  g0965(.a(n1092), .b(n469), .O(n1093));
  orx   g0966(.a(n1093), .b(n471), .O(n1094));
  invx  g0967(.a(n506), .O(n1095));
  andx  g0968(.a(n1095), .b(n1094), .O(n1096));
  andx  g0969(.a(n1096), .b(n499), .O(n1097));
  orx   g0970(.a(n1097), .b(n501), .O(n1098));
  invx  g0971(.a(n536), .O(n1099));
  andx  g0972(.a(n1099), .b(n1098), .O(n1100));
  andx  g0973(.a(n1100), .b(n529), .O(n1101));
  orx   g0974(.a(n1101), .b(n531), .O(n1102));
  invx  g0975(.a(n566), .O(n1103));
  andx  g0976(.a(n1103), .b(n1102), .O(n1104));
  andx  g0977(.a(n1104), .b(n559), .O(n1105));
  orx   g0978(.a(n1105), .b(n561), .O(n1106));
  invx  g0979(.a(n596), .O(n1107));
  andx  g0980(.a(n1107), .b(n1106), .O(n1108));
  andx  g0981(.a(n1108), .b(n589), .O(n1109));
  orx   g0982(.a(n1109), .b(n591), .O(n1110));
  invx  g0983(.a(n626), .O(n1111));
  andx  g0984(.a(n1111), .b(n1110), .O(n1112));
  andx  g0985(.a(n1112), .b(n619), .O(n1113));
  orx   g0986(.a(n1113), .b(n621), .O(n1114));
  invx  g0987(.a(n656), .O(n1115));
  andx  g0988(.a(n1115), .b(n1114), .O(n1116));
  andx  g0989(.a(n1116), .b(n649), .O(n1117));
  orx   g0990(.a(n1117), .b(n651), .O(n1118));
  invx  g0991(.a(n686), .O(n1119));
  andx  g0992(.a(n1119), .b(n1118), .O(n1120));
  andx  g0993(.a(n1120), .b(n679), .O(n1121));
  orx   g0994(.a(n1121), .b(n681), .O(n1122));
  invx  g0995(.a(n716), .O(n1123));
  andx  g0996(.a(n1123), .b(n1122), .O(n1124));
  andx  g0997(.a(n1124), .b(n709), .O(n1125));
  orx   g0998(.a(n1125), .b(n711), .O(n1126));
  invx  g0999(.a(n746), .O(n1127));
  andx  g1000(.a(n1127), .b(n1126), .O(n1128));
  andx  g1001(.a(n1128), .b(n739), .O(n1129));
  orx   g1002(.a(n1129), .b(n741), .O(n1130));
  invx  g1003(.a(n776), .O(n1131));
  andx  g1004(.a(n1131), .b(n1130), .O(n1132));
  andx  g1005(.a(n1132), .b(n769), .O(n1133));
  orx   g1006(.a(n1133), .b(n771), .O(n1134));
  invx  g1007(.a(n806), .O(n1135));
  andx  g1008(.a(n1135), .b(n1134), .O(n1136));
  andx  g1009(.a(n1136), .b(n799), .O(n1137));
  orx   g1010(.a(n1137), .b(n801), .O(n1138));
  invx  g1011(.a(n836), .O(n1139));
  andx  g1012(.a(n1139), .b(n1138), .O(n1140));
  andx  g1013(.a(n1140), .b(n829), .O(n1141));
  orx   g1014(.a(n1141), .b(n831), .O(n1142));
  invx  g1015(.a(n866), .O(n1143));
  andx  g1016(.a(n1143), .b(n1142), .O(n1144));
  andx  g1017(.a(n1144), .b(n859), .O(n1145));
  orx   g1018(.a(n1145), .b(n861), .O(n1146));
  invx  g1019(.a(n896), .O(n1147));
  andx  g1020(.a(n1147), .b(n1146), .O(n1148));
  andx  g1021(.a(n1148), .b(n889), .O(n1149));
  orx   g1022(.a(n1149), .b(n891), .O(n1150));
  invx  g1023(.a(n926), .O(n1151));
  andx  g1024(.a(n1151), .b(n1150), .O(n1152));
  andx  g1025(.a(n1152), .b(n919), .O(n1153));
  orx   g1026(.a(n1153), .b(n921), .O(n1154));
  invx  g1027(.a(n956), .O(n1155));
  andx  g1028(.a(n1155), .b(n1154), .O(n1156));
  andx  g1029(.a(n1156), .b(n949), .O(n1157));
  orx   g1030(.a(n1157), .b(n951), .O(n1158));
  invx  g1031(.a(n986), .O(n1159));
  andx  g1032(.a(n1159), .b(n1158), .O(n1160));
  andx  g1033(.a(n1160), .b(n979), .O(n1161));
  orx   g1034(.a(n1161), .b(n981), .O(n1162));
  invx  g1035(.a(n1016), .O(n1163));
  andx  g1036(.a(n1163), .b(n1162), .O(n1164));
  andx  g1037(.a(n1164), .b(n1009), .O(n1165));
  orx   g1038(.a(n1165), .b(n1011), .O(n1166));
  invx  g1039(.a(n1047), .O(n1167));
  andx  g1040(.a(n1167), .b(n1166), .O(n1168));
  orx   g1041(.a(n1168), .b(n1043), .O(n1169));
  andx  g1042(.a(n1169), .b(n1049), .O(n1170));
  andx  g1043(.a(n1170), .b(pi95), .O(n1171));
  invx  g1044(.a(pi95), .O(n1172));
  andx  g1045(.a(n1168), .b(n1043), .O(n1173));
  andx  g1046(.a(n1048), .b(n1044), .O(n1174));
  orx   g1047(.a(n1174), .b(n1173), .O(n1175));
  andx  g1048(.a(n1175), .b(n1172), .O(n1176));
  orx   g1049(.a(n1176), .b(n1171), .O(n1177));
  orx   g1050(.a(n1030), .b(n1021), .O(n1178));
  andx  g1051(.a(n1178), .b(pi92), .O(n1179));
  andx  g1052(.a(n1030), .b(n1021), .O(n1180));
  orx   g1053(.a(n1180), .b(n1179), .O(n1181));
  andx  g1054(.a(n1181), .b(n1177), .O(n1182));
  orx   g1055(.a(n1175), .b(n1172), .O(n1183));
  orx   g1056(.a(n1170), .b(pi95), .O(n1184));
  andx  g1057(.a(n1184), .b(n1183), .O(n1185));
  andx  g1058(.a(n1036), .b(n1024), .O(n1186));
  orx   g1059(.a(n1186), .b(n1023), .O(n1187));
  orx   g1060(.a(n1036), .b(n1024), .O(n1188));
  andx  g1061(.a(n1188), .b(n1187), .O(n1189));
  andx  g1062(.a(n1189), .b(n1185), .O(n1190));
  orx   g1063(.a(n1190), .b(n1182), .O(po31));
endmodule


