// Benchmark "top" written by ABC on Fri Feb  7 13:33:15 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25;
  wire n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n97, n99, n100,
    n101, n103, n105, n106, n107, n108, n109, n110, n111, n114, n115, n116,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n189, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n283, n285, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n366, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n384, n386, n387, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n408, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447;
  xorx g000(.a(pi38), .b(pi45), .O(n86));
  xorx g001(.a(n86), .b(pi02), .O(n87));
  invx g002(.a(pi01), .O(n88));
  xorx g003(.a(pi21), .b(pi25), .O(n89));
  xorx g004(.a(n89), .b(n88), .O(n90));
  xorx g005(.a(n90), .b(n87), .O(n91));
  xorx g006(.a(pi15), .b(pi19), .O(n92));
  invx g007(.a(pi47), .O(n93));
  xorx g008(.a(pi48), .b(n93), .O(n94));
  xorx g009(.a(n94), .b(n92), .O(n95));
  xorx g010(.a(n95), .b(n91), .O(po00));
  andx g011(.a(pi28), .b(pi30), .O(n97));
  andx g012(.a(n97), .b(pi13), .O(po01));
  invx g013(.a(pi31), .O(n99));
  andx g014(.a(pi12), .b(pi28), .O(n100));
  invx g015(.a(n100), .O(n101));
  orx  g016(.a(n101), .b(n99), .O(po02));
  orx  g017(.a(pi54), .b(pi55), .O(n103));
  andx g018(.a(n103), .b(pi56), .O(po03));
  andx g019(.a(pi35), .b(pi07), .O(n105));
  invx g020(.a(n105), .O(n106));
  invx g021(.a(pi29), .O(n107));
  invx g022(.a(pi33), .O(n108));
  orx  g023(.a(n108), .b(n107), .O(n109));
  orx  g024(.a(n109), .b(n106), .O(n110));
  andx g025(.a(pi08), .b(pi30), .O(n111));
  andx g026(.a(n111), .b(pi13), .O(po24));
  orx  g027(.a(po24), .b(n110), .O(po04));
  invx g028(.a(pi48), .O(n114));
  invx g029(.a(pi46), .O(n115));
  andx g030(.a(pi34), .b(pi35), .O(n116));
  andx g031(.a(n116), .b(pi33), .O(po14));
  andx g032(.a(pi32), .b(pi31), .O(n118));
  xorx g033(.a(pi29), .b(pi30), .O(n119));
  andx g034(.a(n119), .b(n118), .O(n120));
  andx g035(.a(n120), .b(po14), .O(n121));
  invx g036(.a(n121), .O(n122));
  andx g037(.a(n97), .b(pi31), .O(n123));
  andx g038(.a(pi26), .b(pi29), .O(n124));
  andx g039(.a(n124), .b(n116), .O(n125));
  invx g040(.a(n125), .O(n126));
  orx  g041(.a(n126), .b(n123), .O(n127));
  andx g042(.a(n127), .b(n122), .O(n128));
  orx  g043(.a(n128), .b(n115), .O(n129));
  andx g044(.a(n100), .b(pi13), .O(n130));
  andx g045(.a(n130), .b(po14), .O(n131));
  invx g046(.a(pi14), .O(n132));
  andx g047(.a(n132), .b(pi27), .O(n133));
  andx g048(.a(n133), .b(n131), .O(n134));
  invx g049(.a(n134), .O(n135));
  invx g050(.a(pi41), .O(n136));
  invx g051(.a(pi35), .O(n137));
  invx g052(.a(pi34), .O(n138));
  orx  g053(.a(n138), .b(n137), .O(n139));
  orx  g054(.a(n139), .b(n108), .O(n140));
  orx  g055(.a(n118), .b(n107), .O(n141));
  orx  g056(.a(n141), .b(n140), .O(n142));
  andx g057(.a(n142), .b(pi35), .O(n143));
  orx  g058(.a(n143), .b(n136), .O(n144));
  andx g059(.a(n144), .b(n135), .O(n145));
  andx g060(.a(n145), .b(n129), .O(n146));
  orx  g061(.a(n146), .b(n114), .O(n147));
  invx g062(.a(n123), .O(n148));
  andx g063(.a(n125), .b(n148), .O(n149));
  orx  g064(.a(n149), .b(n121), .O(n150));
  andx g065(.a(n150), .b(pi46), .O(n151));
  invx g066(.a(pi32), .O(n152));
  orx  g067(.a(n152), .b(n99), .O(n153));
  andx g068(.a(n153), .b(pi29), .O(n154));
  andx g069(.a(n154), .b(po14), .O(n155));
  orx  g070(.a(n155), .b(n137), .O(n156));
  andx g071(.a(n156), .b(pi41), .O(n157));
  orx  g072(.a(n157), .b(n134), .O(n158));
  orx  g073(.a(n158), .b(n151), .O(n159));
  orx  g074(.a(n159), .b(pi48), .O(n160));
  andx g075(.a(n160), .b(n147), .O(n161));
  orx  g076(.a(n161), .b(pi49), .O(n162));
  andx g077(.a(n159), .b(pi48), .O(n163));
  invx g078(.a(pi49), .O(n164));
  andx g079(.a(n146), .b(n114), .O(n165));
  orx  g080(.a(n165), .b(n164), .O(n166));
  orx  g081(.a(n166), .b(n163), .O(n167));
  andx g082(.a(n167), .b(pi36), .O(n168));
  andx g083(.a(n168), .b(n162), .O(n169));
  andx g084(.a(n161), .b(pi11), .O(n170));
  andx g085(.a(n163), .b(pi09), .O(n171));
  andx g086(.a(n159), .b(pi10), .O(n172));
  andx g087(.a(pi27), .b(pi26), .O(n173));
  andx g088(.a(n173), .b(n105), .O(n174));
  andx g089(.a(pi05), .b(pi31), .O(n175));
  andx g090(.a(pi03), .b(pi30), .O(n176));
  andx g091(.a(n176), .b(pi04), .O(n177));
  andx g092(.a(n177), .b(n175), .O(n178));
  andx g093(.a(n178), .b(n174), .O(n179));
  andx g094(.a(n179), .b(pi48), .O(n180));
  andx g095(.a(pi53), .b(pi51), .O(n181));
  andx g096(.a(pi16), .b(pi43), .O(n182));
  orx  g097(.a(n182), .b(n181), .O(n183));
  orx  g098(.a(n183), .b(n180), .O(n184));
  orx  g099(.a(n184), .b(n172), .O(n185));
  orx  g100(.a(n185), .b(n171), .O(n186));
  orx  g101(.a(n186), .b(n170), .O(n187));
  orx  g102(.a(n187), .b(n169), .O(po05));
  andx g103(.a(pi08), .b(pi12), .O(n189));
  andx g104(.a(n189), .b(pi13), .O(po06));
  xorx g105(.a(pi40), .b(pi39), .O(n191));
  xorx g106(.a(n191), .b(pi00), .O(n192));
  xorx g107(.a(pi20), .b(pi22), .O(n193));
  xorx g108(.a(n193), .b(n88), .O(n194));
  xorx g109(.a(n194), .b(n192), .O(n195));
  xorx g110(.a(pi17), .b(pi18), .O(n196));
  invx g111(.a(pi43), .O(n197));
  xorx g112(.a(pi46), .b(n197), .O(n198));
  xorx g113(.a(n198), .b(n196), .O(n199));
  xorx g114(.a(n199), .b(n195), .O(po07));
  andx g115(.a(n150), .b(pi22), .O(n201));
  andx g116(.a(n132), .b(pi29), .O(n202));
  andx g117(.a(n202), .b(n131), .O(n203));
  andx g118(.a(pi23), .b(pi24), .O(n204));
  andx g119(.a(n153), .b(pi27), .O(n205));
  andx g120(.a(n205), .b(po14), .O(n206));
  andx g121(.a(n206), .b(pi41), .O(n207));
  orx  g122(.a(n207), .b(n204), .O(n208));
  orx  g123(.a(n208), .b(n203), .O(n209));
  orx  g124(.a(n209), .b(n201), .O(n210));
  andx g125(.a(n210), .b(pi25), .O(n211));
  invx g126(.a(n211), .O(n212));
  orx  g127(.a(n210), .b(pi25), .O(n213));
  andx g128(.a(n213), .b(n212), .O(n214));
  invx g129(.a(n214), .O(n215));
  andx g130(.a(n166), .b(n147), .O(n216));
  invx g131(.a(pi45), .O(n217));
  andx g132(.a(n150), .b(pi40), .O(n218));
  invx g133(.a(n218), .O(n219));
  invx g134(.a(pi42), .O(n220));
  orx  g135(.a(n143), .b(n220), .O(n221));
  andx g136(.a(n221), .b(n135), .O(n222));
  andx g137(.a(n222), .b(n219), .O(n223));
  andx g138(.a(n223), .b(n217), .O(n224));
  andx g139(.a(n150), .b(pi43), .O(n225));
  invx g140(.a(n225), .O(n226));
  invx g141(.a(pi44), .O(n227));
  orx  g142(.a(n143), .b(n227), .O(n228));
  andx g143(.a(n228), .b(n135), .O(n229));
  andx g144(.a(n229), .b(n226), .O(n230));
  andx g145(.a(n230), .b(n93), .O(n231));
  orx  g146(.a(n231), .b(n224), .O(n232));
  orx  g147(.a(n232), .b(n216), .O(n233));
  orx  g148(.a(n230), .b(n93), .O(n234));
  orx  g149(.a(n234), .b(n224), .O(n235));
  andx g150(.a(n156), .b(pi42), .O(n236));
  orx  g151(.a(n236), .b(n134), .O(n237));
  orx  g152(.a(n237), .b(n218), .O(n238));
  andx g153(.a(n238), .b(pi45), .O(n239));
  invx g154(.a(n239), .O(n240));
  andx g155(.a(n240), .b(n235), .O(n241));
  andx g156(.a(n241), .b(n233), .O(n242));
  andx g157(.a(n150), .b(pi39), .O(n243));
  andx g158(.a(n156), .b(pi37), .O(n244));
  orx  g159(.a(n244), .b(n134), .O(n245));
  orx  g160(.a(n245), .b(n243), .O(n246));
  orx  g161(.a(n246), .b(pi38), .O(n247));
  invx g162(.a(n247), .O(n248));
  orx  g163(.a(n248), .b(n242), .O(n249));
  andx g164(.a(n246), .b(pi38), .O(n250));
  invx g165(.a(n250), .O(n251));
  andx g166(.a(n251), .b(n249), .O(n252));
  orx  g167(.a(n252), .b(n215), .O(n253));
  andx g168(.a(n160), .b(pi49), .O(n254));
  orx  g169(.a(n254), .b(n163), .O(n255));
  orx  g170(.a(n238), .b(pi45), .O(n256));
  andx g171(.a(n156), .b(pi44), .O(n257));
  orx  g172(.a(n257), .b(n134), .O(n258));
  orx  g173(.a(n258), .b(n225), .O(n259));
  orx  g174(.a(n259), .b(pi47), .O(n260));
  andx g175(.a(n260), .b(n256), .O(n261));
  andx g176(.a(n261), .b(n255), .O(n262));
  andx g177(.a(n259), .b(pi47), .O(n263));
  andx g178(.a(n263), .b(n256), .O(n264));
  orx  g179(.a(n239), .b(n264), .O(n265));
  orx  g180(.a(n265), .b(n262), .O(n266));
  andx g181(.a(n247), .b(n266), .O(n267));
  orx  g182(.a(n250), .b(n267), .O(n268));
  orx  g183(.a(n268), .b(n214), .O(n269));
  andx g184(.a(n269), .b(pi36), .O(n270));
  andx g185(.a(n270), .b(n253), .O(n271));
  andx g186(.a(n214), .b(pi11), .O(n272));
  andx g187(.a(n211), .b(pi09), .O(n273));
  andx g188(.a(n210), .b(pi10), .O(n274));
  andx g189(.a(n179), .b(pi25), .O(n275));
  andx g190(.a(pi20), .b(pi16), .O(n276));
  orx  g191(.a(n276), .b(n275), .O(n277));
  orx  g192(.a(n277), .b(n274), .O(n278));
  orx  g193(.a(n278), .b(n273), .O(n279));
  orx  g194(.a(n279), .b(n272), .O(n280));
  orx  g195(.a(n280), .b(n271), .O(po08));
  andx g196(.a(n124), .b(n105), .O(po09));
  invx g197(.a(n189), .O(n283));
  orx  g198(.a(n283), .b(n99), .O(po10));
  invx g199(.a(n111), .O(n285));
  orx  g200(.a(n285), .b(n99), .O(po11));
  andx g201(.a(n150), .b(pi17), .O(n287));
  andx g202(.a(pi24), .b(pi26), .O(n288));
  andx g203(.a(n206), .b(pi37), .O(n289));
  orx  g204(.a(n289), .b(n288), .O(n290));
  orx  g205(.a(n290), .b(n203), .O(n291));
  orx  g206(.a(n291), .b(n287), .O(n292));
  xorx g207(.a(n292), .b(pi15), .O(n293));
  invx g208(.a(n293), .O(n294));
  invx g209(.a(n213), .O(n295));
  orx  g210(.a(n252), .b(n295), .O(n296));
  andx g211(.a(n150), .b(pi20), .O(n297));
  andx g212(.a(pi24), .b(pi29), .O(n298));
  andx g213(.a(n206), .b(pi44), .O(n299));
  orx  g214(.a(n299), .b(n298), .O(n300));
  orx  g215(.a(n300), .b(n203), .O(n301));
  orx  g216(.a(n301), .b(n297), .O(n302));
  orx  g217(.a(n302), .b(pi21), .O(n303));
  invx g218(.a(pi19), .O(n304));
  andx g219(.a(n150), .b(pi18), .O(n305));
  andx g220(.a(pi24), .b(pi34), .O(n306));
  andx g221(.a(n206), .b(pi42), .O(n307));
  orx  g222(.a(n307), .b(n306), .O(n308));
  orx  g223(.a(n308), .b(n203), .O(n309));
  orx  g224(.a(n309), .b(n305), .O(n310));
  invx g225(.a(n310), .O(n311));
  andx g226(.a(n311), .b(n304), .O(n312));
  invx g227(.a(n312), .O(n313));
  andx g228(.a(n313), .b(n303), .O(n314));
  invx g229(.a(n314), .O(n315));
  orx  g230(.a(n315), .b(n296), .O(n316));
  andx g231(.a(n302), .b(pi21), .O(n317));
  orx  g232(.a(n317), .b(n211), .O(n318));
  andx g233(.a(n318), .b(n303), .O(n319));
  andx g234(.a(n319), .b(n313), .O(n320));
  andx g235(.a(n310), .b(pi19), .O(n321));
  orx  g236(.a(n321), .b(n320), .O(n322));
  invx g237(.a(n322), .O(n323));
  andx g238(.a(n323), .b(n316), .O(n324));
  orx  g239(.a(n324), .b(n294), .O(n325));
  andx g240(.a(n268), .b(n213), .O(n326));
  andx g241(.a(n314), .b(n326), .O(n327));
  orx  g242(.a(n322), .b(n327), .O(n328));
  orx  g243(.a(n328), .b(n293), .O(n329));
  andx g244(.a(n329), .b(pi36), .O(n330));
  andx g245(.a(n330), .b(n325), .O(n331));
  andx g246(.a(n293), .b(pi11), .O(n332));
  andx g247(.a(n292), .b(pi15), .O(n333));
  andx g248(.a(n333), .b(pi09), .O(n334));
  andx g249(.a(n292), .b(pi10), .O(n335));
  andx g250(.a(n179), .b(pi15), .O(n336));
  andx g251(.a(pi14), .b(pi16), .O(n337));
  orx  g252(.a(n337), .b(n336), .O(n338));
  orx  g253(.a(n338), .b(n335), .O(n339));
  orx  g254(.a(n339), .b(n334), .O(n340));
  orx  g255(.a(n340), .b(n332), .O(n341));
  orx  g256(.a(n341), .b(n331), .O(po12));
  andx g257(.a(n103), .b(pi57), .O(po13));
  orx  g258(.a(n321), .b(n312), .O(n344));
  invx g259(.a(n344), .O(n345));
  andx g260(.a(n303), .b(n326), .O(n346));
  orx  g261(.a(n346), .b(n319), .O(n347));
  orx  g262(.a(n347), .b(n345), .O(n348));
  invx g263(.a(n319), .O(n349));
  invx g264(.a(n303), .O(n350));
  orx  g265(.a(n350), .b(n296), .O(n351));
  andx g266(.a(n351), .b(n349), .O(n352));
  orx  g267(.a(n352), .b(n344), .O(n353));
  andx g268(.a(n353), .b(pi36), .O(n354));
  andx g269(.a(n354), .b(n348), .O(n355));
  andx g270(.a(n345), .b(pi11), .O(n356));
  andx g271(.a(n321), .b(pi09), .O(n357));
  andx g272(.a(n310), .b(pi10), .O(n358));
  andx g273(.a(n179), .b(pi19), .O(n359));
  andx g274(.a(pi17), .b(pi16), .O(n360));
  orx  g275(.a(n360), .b(n359), .O(n361));
  orx  g276(.a(n361), .b(n358), .O(n362));
  orx  g277(.a(n362), .b(n357), .O(n363));
  orx  g278(.a(n363), .b(n356), .O(n364));
  orx  g279(.a(n364), .b(n355), .O(po15));
  andx g280(.a(n175), .b(pi06), .O(n366));
  andx g281(.a(n366), .b(n174), .O(po16));
  andx g282(.a(n251), .b(n247), .O(n368));
  invx g283(.a(n368), .O(n369));
  orx  g284(.a(n369), .b(n242), .O(n370));
  orx  g285(.a(n368), .b(n266), .O(n371));
  andx g286(.a(n371), .b(pi36), .O(n372));
  andx g287(.a(n372), .b(n370), .O(n373));
  andx g288(.a(n368), .b(pi11), .O(n374));
  andx g289(.a(n250), .b(pi09), .O(n375));
  andx g290(.a(n246), .b(pi10), .O(n376));
  andx g291(.a(n179), .b(pi38), .O(n377));
  andx g292(.a(pi22), .b(pi16), .O(n378));
  orx  g293(.a(n378), .b(n377), .O(n379));
  orx  g294(.a(n379), .b(n376), .O(n380));
  orx  g295(.a(n380), .b(n375), .O(n381));
  orx  g296(.a(n381), .b(n374), .O(n382));
  orx  g297(.a(n382), .b(n373), .O(po17));
  invx g298(.a(po24), .O(n384));
  orx  g299(.a(n384), .b(n110), .O(po18));
  orx  g300(.a(n292), .b(pi15), .O(n386));
  andx g301(.a(n386), .b(n328), .O(n387));
  orx  g302(.a(n387), .b(n333), .O(po19));
  orx  g303(.a(n317), .b(n350), .O(n389));
  invx g304(.a(n389), .O(n390));
  andx g305(.a(n296), .b(n212), .O(n391));
  invx g306(.a(n391), .O(n392));
  orx  g307(.a(n392), .b(n390), .O(n393));
  orx  g308(.a(n391), .b(n389), .O(n394));
  andx g309(.a(n394), .b(pi36), .O(n395));
  andx g310(.a(n395), .b(n393), .O(n396));
  andx g311(.a(n390), .b(pi11), .O(n397));
  andx g312(.a(n317), .b(pi09), .O(n398));
  andx g313(.a(n302), .b(pi10), .O(n399));
  andx g314(.a(n179), .b(pi21), .O(n400));
  andx g315(.a(pi18), .b(pi16), .O(n401));
  orx  g316(.a(n401), .b(n400), .O(n402));
  orx  g317(.a(n402), .b(n399), .O(n403));
  orx  g318(.a(n403), .b(n398), .O(n404));
  orx  g319(.a(n404), .b(n397), .O(n405));
  orx  g320(.a(n405), .b(n396), .O(po20));
  andx g321(.a(pi58), .b(pi59), .O(po21));
  andx g322(.a(pi05), .b(pi13), .O(n408));
  andx g323(.a(n408), .b(n174), .O(po22));
  andx g324(.a(n234), .b(n260), .O(n410));
  invx g325(.a(n410), .O(n411));
  orx  g326(.a(n411), .b(n216), .O(n412));
  orx  g327(.a(n410), .b(n255), .O(n413));
  andx g328(.a(n413), .b(pi36), .O(n414));
  andx g329(.a(n414), .b(n412), .O(n415));
  andx g330(.a(n410), .b(pi11), .O(n416));
  andx g331(.a(n263), .b(pi09), .O(n417));
  andx g332(.a(n259), .b(pi10), .O(n418));
  andx g333(.a(n179), .b(pi47), .O(n419));
  andx g334(.a(pi52), .b(pi51), .O(n420));
  andx g335(.a(pi40), .b(pi16), .O(n421));
  orx  g336(.a(n421), .b(n420), .O(n422));
  orx  g337(.a(n422), .b(n419), .O(n423));
  orx  g338(.a(n423), .b(n418), .O(n424));
  orx  g339(.a(n424), .b(n417), .O(n425));
  orx  g340(.a(n425), .b(n416), .O(n426));
  orx  g341(.a(n426), .b(n415), .O(po23));
  andx g342(.a(n240), .b(n256), .O(n428));
  andx g343(.a(n260), .b(n255), .O(n429));
  orx  g344(.a(n429), .b(n263), .O(n430));
  orx  g345(.a(n430), .b(n428), .O(n431));
  invx g346(.a(n428), .O(n432));
  invx g347(.a(n430), .O(n433));
  orx  g348(.a(n433), .b(n432), .O(n434));
  andx g349(.a(n434), .b(pi36), .O(n435));
  andx g350(.a(n435), .b(n431), .O(n436));
  andx g351(.a(n428), .b(pi11), .O(n437));
  andx g352(.a(n239), .b(pi09), .O(n438));
  andx g353(.a(n238), .b(pi10), .O(n439));
  andx g354(.a(n179), .b(pi45), .O(n440));
  andx g355(.a(pi50), .b(pi51), .O(n441));
  andx g356(.a(pi39), .b(pi16), .O(n442));
  orx  g357(.a(n442), .b(n441), .O(n443));
  orx  g358(.a(n443), .b(n440), .O(n444));
  orx  g359(.a(n444), .b(n439), .O(n445));
  orx  g360(.a(n445), .b(n438), .O(n446));
  orx  g361(.a(n446), .b(n437), .O(n447));
  orx  g362(.a(n447), .b(n436), .O(po25));
endmodule


