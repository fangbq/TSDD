// Benchmark "logsig_approx" written by ABC on Fri Feb  7 13:42:21 2014

module logsig_approx ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29;
  wire n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
    n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
    n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n155, n156, n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n237,
    n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280, n281, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n504, n505, n507, n508, n509, n510, n512, n513, n514,
    n515, n516, n517, n518, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
    n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378;
  bufx g0000(.A(pi22), .O(n62));
  bufx g0001(.A(n1251), .O(n63));
  bufx g0002(.A(n1257), .O(n64));
  bufx g0003(.A(n1248), .O(n65));
  bufx g0004(.A(n1308), .O(n66));
  bufx g0005(.A(n1205), .O(n67));
  bufx g0006(.A(n1271), .O(n68));
  bufx g0007(.A(n1327), .O(n69));
  bufx g0008(.A(n1311), .O(n70));
  bufx g0009(.A(n999), .O(n71));
  bufx g0010(.A(n1286), .O(n72));
  bufx g0011(.A(n1276), .O(n73));
  bufx g0012(.A(n1088), .O(n74));
  bufx g0013(.A(n866), .O(n75));
  bufx g0014(.A(n979), .O(n76));
  bufx g0015(.A(n1028), .O(n77));
  bufx g0016(.A(n1350), .O(n78));
  bufx g0017(.A(n1303), .O(n79));
  bufx g0018(.A(n1215), .O(n80));
  invx g0019(.A(n1252), .O(n81));
  invx g0020(.A(n81), .O(n82));
  bufx g0021(.A(n1318), .O(n83));
  invx g0022(.A(n1203), .O(n84));
  bufx g0023(.A(n1033), .O(n85));
  bufx g0024(.A(n1138), .O(n86));
  invx g0025(.A(n1331), .O(n87));
  invx g0026(.A(n87), .O(n88));
  invx g0027(.A(n1153), .O(n89));
  invx g0028(.A(n89), .O(n90));
  bufx g0029(.A(n1289), .O(n91));
  bufx g0030(.A(n1347), .O(n92));
  invx g0031(.A(n1267), .O(n93));
  invx g0032(.A(n93), .O(n94));
  bufx g0033(.A(n1229), .O(n95));
  invx g0034(.A(n1304), .O(n96));
  invx g0035(.A(n96), .O(n97));
  bufx g0036(.A(n1077), .O(n98));
  bufx g0037(.A(n1279), .O(n99));
  bufx g0038(.A(n1188), .O(n100));
  bufx g0039(.A(n1102), .O(n101));
  bufx g0040(.A(n1059), .O(n102));
  bufx g0041(.A(n1036), .O(n103));
  bufx g0042(.A(n1361), .O(n104));
  bufx g0043(.A(n1237), .O(n105));
  bufx g0044(.A(n1038), .O(n106));
  bufx g0045(.A(n1334), .O(n107));
  bufx g0046(.A(n1297), .O(n108));
  bufx g0047(.A(n1260), .O(n109));
  bufx g0048(.A(n1195), .O(n110));
  invx g0049(.A(n1278), .O(n111));
  invx g0050(.A(n111), .O(n112));
  bufx g0051(.A(n1346), .O(n113));
  bufx g0052(.A(n1346), .O(n114));
  bufx g0053(.A(n960), .O(n115));
  bufx g0054(.A(n1187), .O(n116));
  invx g0055(.A(n373), .O(n117));
  bufx g0056(.A(n1288), .O(n118));
  bufx g0057(.A(n1144), .O(n119));
  bufx g0058(.A(n1177), .O(n120));
  invx g0059(.A(n1362), .O(n121));
  invx g0060(.A(n121), .O(n122));
  invx g0061(.A(n1305), .O(n123));
  invx g0062(.A(n123), .O(n124));
  invx g0063(.A(n1272), .O(n125));
  invx g0064(.A(n125), .O(n126));
  bufx g0065(.A(n1275), .O(n127));
  bufx g0066(.A(n1275), .O(n128));
  bufx g0067(.A(n1307), .O(n129));
  bufx g0068(.A(n1307), .O(n130));
  invx g0069(.A(n1317), .O(n131));
  invx g0070(.A(n131), .O(n132));
  invx g0071(.A(n131), .O(n133));
  bufx g0072(.A(n1265), .O(n134));
  bufx g0073(.A(n504), .O(n135));
  bufx g0074(.A(n1228), .O(n136));
  bufx g0075(.A(n1176), .O(n137));
  bufx g0076(.A(n1326), .O(n138));
  invx g0077(.A(n1315), .O(n139));
  invx g0078(.A(n139), .O(n140));
  invx g0079(.A(n1274), .O(n141));
  invx g0080(.A(n141), .O(n142));
  invx g0081(.A(n141), .O(n143));
  invx g0082(.A(n1363), .O(n144));
  invx g0083(.A(n144), .O(n145));
  invx g0084(.A(n144), .O(n146));
  invx g0085(.A(n1306), .O(n147));
  invx g0086(.A(n147), .O(n148));
  invx g0087(.A(n147), .O(n149));
  bufx g0088(.A(n1364), .O(n150));
  bufx g0089(.A(n1364), .O(n151));
  bufx g0090(.A(n1364), .O(n152));
  bufx g0091(.A(n1364), .O(n153));
  andx g0092(.A(n155), .B(n151), .O(po09));
  orx  g0093(.A(n189), .B(n156), .O(n155));
  andx g0094(.A(n235), .B(n157), .O(n156));
  orx  g0095(.A(n158), .B(n1049), .O(n157));
  andx g0096(.A(n332), .B(n159), .O(n158));
  orx  g0097(.A(n160), .B(n382), .O(n159));
  andx g0098(.A(n373), .B(n161), .O(n160));
  orx  g0099(.A(n162), .B(n926), .O(n161));
  andx g0100(.A(n163), .B(n1038), .O(n162));
  andx g0101(.A(n164), .B(n1182), .O(n163));
  orx  g0102(.A(n165), .B(n116), .O(n164));
  andx g0103(.A(n1035), .B(n166), .O(n165));
  orx  g0104(.A(n167), .B(n98), .O(n166));
  andx g0105(.A(n1310), .B(n168), .O(n167));
  orx  g0106(.A(n169), .B(n110), .O(n168));
  andx g0107(.A(n1130), .B(n170), .O(n169));
  orx  g0108(.A(n171), .B(n1083), .O(n170));
  andx g0109(.A(n966), .B(n172), .O(n171));
  orx  g0110(.A(n173), .B(n108), .O(n172));
  andx g0111(.A(n174), .B(n123), .O(n173));
  orx  g0112(.A(n175), .B(n67), .O(n174));
  andx g0113(.A(n830), .B(n176), .O(n175));
  orx  g0114(.A(n177), .B(n118), .O(n176));
  andx g0115(.A(n178), .B(n147), .O(n177));
  orx  g0116(.A(n179), .B(n400), .O(n178));
  andx g0117(.A(n111), .B(n180), .O(n179));
  orx  g0118(.A(n181), .B(n95), .O(n180));
  andx g0119(.A(n182), .B(n66), .O(n181));
  orx  g0120(.A(n183), .B(n896), .O(n182));
  andx g0121(.A(n184), .B(n1242), .O(n183));
  orx  g0122(.A(n185), .B(n63), .O(n184));
  andx g0123(.A(n413), .B(n186), .O(n185));
  orx  g0124(.A(n187), .B(n1266), .O(n186));
  andx g0125(.A(n904), .B(n188), .O(n187));
  orx  g0126(.A(pi09), .B(n757), .O(n188));
  andx g0127(.A(n1353), .B(n1041), .O(n189));
  andx g0128(.A(n191), .B(n150), .O(po08));
  orx  g0129(.A(n192), .B(n548), .O(n191));
  andx g0130(.A(n235), .B(n193), .O(n192));
  orx  g0131(.A(n194), .B(n1362), .O(n193));
  andx g0132(.A(n1146), .B(n195), .O(n194));
  orx  g0133(.A(n196), .B(n330), .O(n195));
  andx g0134(.A(n908), .B(n197), .O(n196));
  orx  g0135(.A(n198), .B(n102), .O(n197));
  andx g0136(.A(n1141), .B(n199), .O(n198));
  orx  g0137(.A(n200), .B(n88), .O(n199));
  andx g0138(.A(n1065), .B(n201), .O(n200));
  orx  g0139(.A(n202), .B(n138), .O(n201));
  andx g0140(.A(n1175), .B(n203), .O(n202));
  orx  g0141(.A(n204), .B(n1173), .O(n203));
  andx g0142(.A(n205), .B(n1365), .O(n204));
  orx  g0143(.A(n206), .B(n1183), .O(n205));
  andx g0144(.A(n207), .B(n139), .O(n206));
  orx  g0145(.A(n208), .B(n86), .O(n207));
  andx g0146(.A(n1035), .B(n209), .O(n208));
  orx  g0147(.A(n210), .B(n1135), .O(n209));
  andx g0148(.A(n1310), .B(n211), .O(n210));
  orx  g0149(.A(n71), .B(n212), .O(n211));
  orx  g0150(.A(n79), .B(n213), .O(n212));
  andx g0151(.A(n758), .B(n214), .O(n213));
  orx  g0152(.A(n215), .B(n303), .O(n214));
  andx g0153(.A(n1292), .B(n216), .O(n215));
  orx  g0154(.A(n217), .B(n694), .O(n216));
  andx g0155(.A(n115), .B(n218), .O(n217));
  orx  g0156(.A(n219), .B(n101), .O(n218));
  andx g0157(.A(n1282), .B(n220), .O(n219));
  orx  g0158(.A(n221), .B(n703), .O(n220));
  andx g0159(.A(n905), .B(n222), .O(n221));
  orx  g0160(.A(n95), .B(n223), .O(n222));
  orx  g0161(.A(n1110), .B(n224), .O(n223));
  andx g0162(.A(n225), .B(n1123), .O(n224));
  andx g0163(.A(n226), .B(n1232), .O(n225));
  orx  g0164(.A(n227), .B(n126), .O(n226));
  andx g0165(.A(n1270), .B(n228), .O(n227));
  orx  g0166(.A(n229), .B(n105), .O(n228));
  andx g0167(.A(n230), .B(n1242), .O(n229));
  orx  g0168(.A(n231), .B(n1245), .O(n230));
  andx g0169(.A(n81), .B(n232), .O(n231));
  orx  g0170(.A(n63), .B(n233), .O(n232));
  orx  g0171(.A(n234), .B(n1262), .O(n233));
  andx g0172(.A(pi08), .B(n73), .O(n234));
  invx g0173(.A(n915), .O(n235));
  andx g0174(.A(n1040), .B(n237), .O(po07));
  orx  g0175(.A(n238), .B(n76), .O(n237));
  andx g0176(.A(n1349), .B(n239), .O(n238));
  orx  g0177(.A(n240), .B(n92), .O(n239));
  andx g0178(.A(n1143), .B(n241), .O(n240));
  orx  g0179(.A(n242), .B(n145), .O(n241));
  andx g0180(.A(n1039), .B(n243), .O(n242));
  orx  g0181(.A(n244), .B(n107), .O(n243));
  andx g0182(.A(n373), .B(n245), .O(n244));
  orx  g0183(.A(n246), .B(n1164), .O(n245));
  andx g0184(.A(n599), .B(n247), .O(n246));
  orx  g0185(.A(n248), .B(n138), .O(n247));
  andx g0186(.A(n106), .B(n249), .O(n248));
  orx  g0187(.A(pi30), .B(n250), .O(n249));
  andx g0188(.A(n251), .B(n1182), .O(n250));
  orx  g0189(.A(n252), .B(n1071), .O(n251));
  andx g0190(.A(n1035), .B(n253), .O(n252));
  orx  g0191(.A(n254), .B(n132), .O(n253));
  andx g0192(.A(n759), .B(n255), .O(n254));
  orx  g0193(.A(n256), .B(n1002), .O(n255));
  andx g0194(.A(n648), .B(n257), .O(n256));
  orx  g0195(.A(n258), .B(n71), .O(n257));
  andx g0196(.A(n966), .B(n259), .O(n258));
  orx  g0197(.A(n260), .B(n108), .O(n259));
  andx g0198(.A(n1203), .B(n261), .O(n260));
  orx  g0199(.A(n262), .B(n118), .O(n261));
  andx g0200(.A(n1034), .B(n263), .O(n262));
  orx  g0201(.A(n264), .B(n101), .O(n263));
  andx g0202(.A(n265), .B(n699), .O(n264));
  orx  g0203(.A(n266), .B(n906), .O(n265));
  andx g0204(.A(n1282), .B(n267), .O(n266));
  orx  g0205(.A(n268), .B(n85), .O(n267));
  andx g0206(.A(n851), .B(n269), .O(n268));
  orx  g0207(.A(n270), .B(n80), .O(n269));
  andx g0208(.A(n1029), .B(n271), .O(n270));
  orx  g0209(.A(n272), .B(n95), .O(n271));
  andx g0210(.A(n281), .B(n273), .O(n272));
  orx  g0211(.A(n274), .B(n1226), .O(n273));
  andx g0212(.A(n1122), .B(n275), .O(n274));
  orx  g0213(.A(n276), .B(n1252), .O(n275));
  andx g0214(.A(n1250), .B(n277), .O(n276));
  orx  g0215(.A(n278), .B(n94), .O(n277));
  andx g0216(.A(n413), .B(n279), .O(n278));
  orx  g0217(.A(n128), .B(n280), .O(n279));
  andx g0218(.A(pi07), .B(n1261), .O(n280));
  andx g0219(.A(n589), .B(n66), .O(n281));
  andx g0220(.A(n1040), .B(n283), .O(po06));
  orx  g0221(.A(n284), .B(n1353), .O(n283));
  andx g0222(.A(n1044), .B(n285), .O(n284));
  orx  g0223(.A(n286), .B(n76), .O(n285));
  andx g0224(.A(n1338), .B(n287), .O(n286));
  orx  g0225(.A(n288), .B(n102), .O(n287));
  andx g0226(.A(n1333), .B(n289), .O(n288));
  orx  g0227(.A(n290), .B(n1160), .O(n289));
  andx g0228(.A(n373), .B(n291), .O(n290));
  orx  g0229(.A(n292), .B(n75), .O(n291));
  andx g0230(.A(n1065), .B(n293), .O(n292));
  orx  g0231(.A(n294), .B(n869), .O(n293));
  andx g0232(.A(n724), .B(n295), .O(n294));
  orx  g0233(.A(n1140), .B(n296), .O(n295));
  orx  g0234(.A(n297), .B(n103), .O(n296));
  andx g0235(.A(n1134), .B(n298), .O(n297));
  orx  g0236(.A(n299), .B(n110), .O(n298));
  andx g0237(.A(n801), .B(n300), .O(n299));
  orx  g0238(.A(n97), .B(n301), .O(n300));
  andx g0239(.A(n1129), .B(n302), .O(n301));
  orx  g0240(.A(n305), .B(n303), .O(n302));
  orx  g0241(.A(n304), .B(n1296), .O(n303));
  andx g0242(.A(n67), .B(n123), .O(n304));
  andx g0243(.A(n1096), .B(n306), .O(n305));
  orx  g0244(.A(n307), .B(n118), .O(n306));
  andx g0245(.A(n1034), .B(n308), .O(n307));
  orx  g0246(.A(n72), .B(n309), .O(n308));
  andx g0247(.A(n790), .B(n310), .O(n309));
  orx  g0248(.A(n311), .B(n85), .O(n310));
  andx g0249(.A(n851), .B(n312), .O(n311));
  orx  g0250(.A(n313), .B(n1030), .O(n312));
  andx g0251(.A(n111), .B(n314), .O(n313));
  orx  g0252(.A(n315), .B(n1125), .O(n314));
  andx g0253(.A(n316), .B(n66), .O(n315));
  orx  g0254(.A(n317), .B(n896), .O(n316));
  andx g0255(.A(n1270), .B(n318), .O(n317));
  orx  g0256(.A(n319), .B(n105), .O(n318));
  andx g0257(.A(n1121), .B(n320), .O(n319));
  orx  g0258(.A(n321), .B(n1252), .O(n320));
  andx g0259(.A(n93), .B(n322), .O(n321));
  orx  g0260(.A(n323), .B(n1266), .O(n322));
  andx g0261(.A(n109), .B(pi06), .O(n323));
  andx g0262(.A(n325), .B(n153), .O(po05));
  orx  g0263(.A(n326), .B(n1353), .O(n325));
  andx g0264(.A(n1044), .B(n327), .O(n326));
  orx  g0265(.A(n328), .B(n915), .O(n327));
  andx g0266(.A(n329), .B(n121), .O(n328));
  orx  g0267(.A(n333), .B(n330), .O(n329));
  orx  g0268(.A(n331), .B(n90), .O(n330));
  andx g0269(.A(n332), .B(n78), .O(n331));
  invx g0270(.A(n76), .O(n332));
  andx g0271(.A(n969), .B(n334), .O(n333));
  orx  g0272(.A(n335), .B(n119), .O(n334));
  andx g0273(.A(n1142), .B(n336), .O(n335));
  orx  g0274(.A(n337), .B(n107), .O(n336));
  andx g0275(.A(n373), .B(n338), .O(n337));
  orx  g0276(.A(n339), .B(n75), .O(n338));
  andx g0277(.A(n599), .B(n340), .O(n339));
  orx  g0278(.A(n341), .B(n138), .O(n340));
  andx g0279(.A(n372), .B(n342), .O(n341));
  orx  g0280(.A(n343), .B(n1170), .O(n342));
  andx g0281(.A(n724), .B(n344), .O(n343));
  orx  g0282(.A(n345), .B(n1140), .O(n344));
  andx g0283(.A(n346), .B(n139), .O(n345));
  orx  g0284(.A(n347), .B(n103), .O(n346));
  andx g0285(.A(n1134), .B(n348), .O(n347));
  orx  g0286(.A(n349), .B(n477), .O(n348));
  andx g0287(.A(n1001), .B(n350), .O(n349));
  orx  g0288(.A(n351), .B(n645), .O(n350));
  andx g0289(.A(n352), .B(n648), .O(n351));
  andx g0290(.A(n353), .B(n1301), .O(n352));
  orx  g0291(.A(n354), .B(n79), .O(n353));
  andx g0292(.A(n355), .B(n96), .O(n354));
  orx  g0293(.A(n356), .B(n688), .O(n355));
  andx g0294(.A(n830), .B(n357), .O(n356));
  orx  g0295(.A(n358), .B(n118), .O(n357));
  andx g0296(.A(n359), .B(n147), .O(n358));
  orx  g0297(.A(n360), .B(n961), .O(n359));
  andx g0298(.A(n790), .B(n361), .O(n360));
  orx  g0299(.A(n362), .B(n80), .O(n361));
  andx g0300(.A(n1029), .B(n363), .O(n362));
  orx  g0301(.A(n364), .B(n112), .O(n363));
  andx g0302(.A(n365), .B(n66), .O(n364));
  orx  g0303(.A(n1226), .B(n366), .O(n365));
  andx g0304(.A(n367), .B(n1242), .O(n366));
  orx  g0305(.A(n82), .B(n368), .O(n367));
  orx  g0306(.A(n369), .B(n1247), .O(n368));
  andx g0307(.A(n134), .B(n370), .O(n369));
  orx  g0308(.A(n1262), .B(n371), .O(n370));
  orx  g0309(.A(pi05), .B(n128), .O(n371));
  invx g0310(.A(n120), .O(n372));
  invx g0311(.A(n987), .O(n373));
  andx g0312(.A(n375), .B(n152), .O(po04));
  orx  g0313(.A(n1359), .B(n376), .O(n375));
  andx g0314(.A(n1352), .B(n377), .O(n376));
  orx  g0315(.A(n378), .B(n976), .O(n377));
  andx g0316(.A(n1349), .B(n379), .O(n378));
  orx  g0317(.A(n380), .B(n119), .O(n379));
  andx g0318(.A(n381), .B(n144), .O(n380));
  orx  g0319(.A(n384), .B(n382), .O(n381));
  orx  g0320(.A(n383), .B(n1339), .O(n382));
  andx g0321(.A(n1039), .B(n107), .O(n383));
  andx g0322(.A(n852), .B(n385), .O(n384));
  orx  g0323(.A(n386), .B(n1164), .O(n385));
  andx g0324(.A(n106), .B(n387), .O(n386));
  orx  g0325(.A(n388), .B(n137), .O(n387));
  andx g0326(.A(n1181), .B(n389), .O(n388));
  orx  g0327(.A(n140), .B(n390), .O(n389));
  andx g0328(.A(n1313), .B(n391), .O(n390));
  orx  g0329(.A(n392), .B(n98), .O(n391));
  andx g0330(.A(n1131), .B(n393), .O(n392));
  orx  g0331(.A(n394), .B(n110), .O(n393));
  andx g0332(.A(n801), .B(n395), .O(n394));
  orx  g0333(.A(n1304), .B(n396), .O(n395));
  andx g0334(.A(n963), .B(n397), .O(n396));
  orx  g0335(.A(n398), .B(n84), .O(n397));
  andx g0336(.A(n115), .B(n399), .O(n398));
  orx  g0337(.A(n402), .B(n400), .O(n399));
  orx  g0338(.A(n401), .B(n581), .O(n400));
  andx g0339(.A(n1282), .B(n661), .O(n401));
  andx g0340(.A(n77), .B(n403), .O(n402));
  orx  g0341(.A(n404), .B(n95), .O(n403));
  andx g0342(.A(n1224), .B(n405), .O(n404));
  orx  g0343(.A(n1272), .B(n406), .O(n405));
  andx g0344(.A(n959), .B(n407), .O(n406));
  orx  g0345(.A(n1274), .B(n408), .O(n407));
  andx g0346(.A(n1121), .B(n409), .O(n408));
  orx  g0347(.A(n410), .B(n94), .O(n409));
  andx g0348(.A(n413), .B(n411), .O(n410));
  orx  g0349(.A(n127), .B(n412), .O(n411));
  andx g0350(.A(pi04), .B(n1261), .O(n412));
  invx g0351(.A(n65), .O(n413));
  andx g0352(.A(n1040), .B(n415), .O(po03));
  orx  g0353(.A(n416), .B(n456), .O(n415));
  andx g0354(.A(n1146), .B(n417), .O(n416));
  orx  g0355(.A(n418), .B(n90), .O(n417));
  andx g0356(.A(n969), .B(n419), .O(n418));
  orx  g0357(.A(n420), .B(n92), .O(n419));
  andx g0358(.A(n1142), .B(n421), .O(n420));
  orx  g0359(.A(n422), .B(n107), .O(n421));
  andx g0360(.A(n1141), .B(n423), .O(n422));
  orx  g0361(.A(n424), .B(n75), .O(n423));
  andx g0362(.A(n1065), .B(n425), .O(n424));
  orx  g0363(.A(n426), .B(n69), .O(n425));
  andx g0364(.A(n106), .B(n427), .O(n426));
  orx  g0365(.A(pi30), .B(n428), .O(n427));
  andx g0366(.A(n803), .B(n429), .O(n428));
  orx  g0367(.A(n430), .B(n86), .O(n429));
  andx g0368(.A(n1130), .B(n431), .O(n430));
  orx  g0369(.A(n432), .B(n83), .O(n431));
  andx g0370(.A(n966), .B(n433), .O(n432));
  orx  g0371(.A(n434), .B(n1304), .O(n433));
  andx g0372(.A(n758), .B(n435), .O(n434));
  orx  g0373(.A(n436), .B(n108), .O(n435));
  andx g0374(.A(n1295), .B(n437), .O(n436));
  orx  g0375(.A(n438), .B(n84), .O(n437));
  andx g0376(.A(n830), .B(n439), .O(n438));
  orx  g0377(.A(n442), .B(n440), .O(n439));
  orx  g0378(.A(n441), .B(n91), .O(n440));
  andx g0379(.A(n1287), .B(n149), .O(n441));
  orx  g0380(.A(n453), .B(n443), .O(n442));
  andx g0381(.A(n905), .B(n444), .O(n443));
  orx  g0382(.A(n445), .B(n1030), .O(n444));
  andx g0383(.A(n111), .B(n446), .O(n445));
  orx  g0384(.A(n447), .B(n95), .O(n446));
  andx g0385(.A(n1224), .B(n448), .O(n447));
  orx  g0386(.A(n449), .B(n623), .O(n448));
  andx g0387(.A(n81), .B(n450), .O(n449));
  orx  g0388(.A(n451), .B(n1266), .O(n450));
  andx g0389(.A(n452), .B(n73), .O(n451));
  orx  g0390(.A(n1262), .B(pi03), .O(n452));
  andx g0391(.A(n1101), .B(n614), .O(n453));
  andx g0392(.A(n455), .B(n151), .O(po02));
  orx  g0393(.A(n458), .B(n456), .O(n455));
  orx  g0394(.A(n1361), .B(n457), .O(n456));
  andx g0395(.A(n1352), .B(n915), .O(n457));
  andx g0396(.A(n459), .B(n121), .O(n458));
  orx  g0397(.A(n78), .B(n460), .O(n459));
  orx  g0398(.A(n462), .B(n461), .O(n460));
  andx g0399(.A(n908), .B(n119), .O(n461));
  andx g0400(.A(n1338), .B(n463), .O(n462));
  orx  g0401(.A(n464), .B(n102), .O(n463));
  andx g0402(.A(n87), .B(n465), .O(n464));
  orx  g0403(.A(n466), .B(n69), .O(n465));
  andx g0404(.A(n1325), .B(n467), .O(n466));
  orx  g0405(.A(n468), .B(n120), .O(n467));
  andx g0406(.A(n106), .B(n469), .O(n468));
  orx  g0407(.A(n470), .B(n721), .O(n469));
  andx g0408(.A(n471), .B(n724), .O(n470));
  andx g0409(.A(n472), .B(n1182), .O(n471));
  orx  g0410(.A(n473), .B(n100), .O(n472));
  andx g0411(.A(n1313), .B(n474), .O(n473));
  orx  g0412(.A(n132), .B(n475), .O(n474));
  andx g0413(.A(n1134), .B(n476), .O(n475));
  orx  g0414(.A(n479), .B(n477), .O(n476));
  orx  g0415(.A(n478), .B(n98), .O(n477));
  andx g0416(.A(n1001), .B(n70), .O(n478));
  andx g0417(.A(n1131), .B(n480), .O(n479));
  orx  g0418(.A(n481), .B(n1081), .O(n480));
  andx g0419(.A(n482), .B(n1130), .O(n481));
  andx g0420(.A(n966), .B(n483), .O(n482));
  orx  g0421(.A(n484), .B(n74), .O(n483));
  andx g0422(.A(n1295), .B(n485), .O(n484));
  orx  g0423(.A(n486), .B(n831), .O(n485));
  andx g0424(.A(n1287), .B(n487), .O(n486));
  orx  g0425(.A(n488), .B(n788), .O(n487));
  andx g0426(.A(n790), .B(n489), .O(n488));
  orx  g0427(.A(n490), .B(n85), .O(n489));
  andx g0428(.A(n77), .B(n491), .O(n490));
  orx  g0429(.A(n1223), .B(n492), .O(n491));
  orx  g0430(.A(n1272), .B(n493), .O(n492));
  andx g0431(.A(n1270), .B(n494), .O(n493));
  orx  g0432(.A(n142), .B(n495), .O(n494));
  andx g0433(.A(n81), .B(n496), .O(n495));
  orx  g0434(.A(n497), .B(n63), .O(n496));
  andx g0435(.A(n109), .B(pi02), .O(n497));
  orx  g0436(.A(pi29), .B(n135), .O(po29));
  orx  g0437(.A(pi28), .B(n135), .O(po28));
  orx  g0438(.A(pi27), .B(n135), .O(po27));
  orx  g0439(.A(pi26), .B(n135), .O(po26));
  orx  g0440(.A(pi25), .B(n135), .O(po25));
  orx  g0441(.A(n505), .B(n135), .O(po24));
  orx  g0442(.A(n1220), .B(n532), .O(n504));
  andx g0443(.A(n1224), .B(pi24), .O(n505));
  orx  g0444(.A(n508), .B(n507), .O(po23));
  invx g0445(.A(n150), .O(n507));
  andx g0446(.A(n509), .B(n1028), .O(n508));
  andx g0447(.A(n801), .B(n510), .O(n509));
  orx  g0448(.A(pi23), .B(n1223), .O(n510));
  andx g0449(.A(n512), .B(n150), .O(po22));
  orx  g0450(.A(n514), .B(n513), .O(n512));
  orx  g0451(.A(n71), .B(n532), .O(n513));
  orx  g0452(.A(n79), .B(n515), .O(n514));
  andx g0453(.A(n77), .B(n516), .O(n515));
  orx  g0454(.A(n1223), .B(n517), .O(n516));
  orx  g0455(.A(n518), .B(n105), .O(n517));
  andx g0456(.A(n81), .B(n62), .O(n518));
  andx g0457(.A(n520), .B(n153), .O(po21));
  orx  g0458(.A(n532), .B(n521), .O(n520));
  orx  g0459(.A(n522), .B(n98), .O(n521));
  andx g0460(.A(n523), .B(n1310), .O(n522));
  andx g0461(.A(n524), .B(n1085), .O(n523));
  orx  g0462(.A(n525), .B(n961), .O(n524));
  andx g0463(.A(n1028), .B(n526), .O(n525));
  orx  g0464(.A(n527), .B(n1223), .O(n526));
  andx g0465(.A(n1122), .B(n528), .O(n527));
  orx  g0466(.A(n529), .B(n63), .O(n528));
  andx g0467(.A(pi21), .B(n73), .O(n529));
  andx g0468(.A(n531), .B(n152), .O(po20));
  orx  g0469(.A(n533), .B(n532), .O(n531));
  orx  g0470(.A(pi30), .B(n1314), .O(n532));
  andx g0471(.A(n759), .B(n534), .O(n533));
  orx  g0472(.A(n535), .B(n110), .O(n534));
  andx g0473(.A(n801), .B(n536), .O(n535));
  orx  g0474(.A(n537), .B(n84), .O(n536));
  andx g0475(.A(n960), .B(n538), .O(n537));
  orx  g0476(.A(n539), .B(n85), .O(n538));
  andx g0477(.A(n1028), .B(n540), .O(n539));
  orx  g0478(.A(n541), .B(n1125), .O(n540));
  andx g0479(.A(n542), .B(n1225), .O(n541));
  orx  g0480(.A(n126), .B(n543), .O(n542));
  andx g0481(.A(n1122), .B(n544), .O(n543));
  orx  g0482(.A(n545), .B(n1244), .O(n544));
  andx g0483(.A(n1250), .B(pi20), .O(n545));
  andx g0484(.A(n547), .B(n151), .O(po01));
  orx  g0485(.A(n551), .B(n548), .O(n547));
  orx  g0486(.A(n549), .B(n1042), .O(n548));
  andx g0487(.A(n1361), .B(n550), .O(n549));
  invx g0488(.A(n1359), .O(n550));
  andx g0489(.A(n89), .B(n552), .O(n551));
  orx  g0490(.A(n553), .B(n76), .O(n552));
  andx g0491(.A(n969), .B(n554), .O(n553));
  orx  g0492(.A(n555), .B(n92), .O(n554));
  andx g0493(.A(n1333), .B(n556), .O(n555));
  orx  g0494(.A(n557), .B(n117), .O(n556));
  andx g0495(.A(n852), .B(n558), .O(n557));
  orx  g0496(.A(n559), .B(n88), .O(n558));
  andx g0497(.A(n599), .B(n560), .O(n559));
  orx  g0498(.A(n561), .B(n138), .O(n560));
  andx g0499(.A(n1175), .B(n562), .O(n561));
  orx  g0500(.A(pi30), .B(n563), .O(n562));
  andx g0501(.A(n564), .B(n1182), .O(n563));
  orx  g0502(.A(n565), .B(n100), .O(n564));
  andx g0503(.A(n566), .B(n139), .O(n565));
  orx  g0504(.A(n567), .B(n86), .O(n566));
  andx g0505(.A(n1035), .B(n568), .O(n567));
  orx  g0506(.A(n569), .B(n1317), .O(n568));
  andx g0507(.A(n1001), .B(n570), .O(n569));
  orx  g0508(.A(n571), .B(n1132), .O(n570));
  andx g0509(.A(n648), .B(n572), .O(n571));
  orx  g0510(.A(n573), .B(n802), .O(n572));
  andx g0511(.A(n574), .B(n96), .O(n573));
  orx  g0512(.A(n575), .B(n883), .O(n574));
  andx g0513(.A(n963), .B(n576), .O(n575));
  orx  g0514(.A(n577), .B(n1206), .O(n576));
  andx g0515(.A(n1128), .B(n578), .O(n577));
  orx  g0516(.A(n579), .B(n828), .O(n578));
  andx g0517(.A(n1287), .B(n580), .O(n579));
  orx  g0518(.A(n583), .B(n581), .O(n580));
  orx  g0519(.A(n582), .B(n101), .O(n581));
  andx g0520(.A(n1282), .B(n99), .O(n582));
  andx g0521(.A(n851), .B(n584), .O(n583));
  orx  g0522(.A(n585), .B(n80), .O(n584));
  andx g0523(.A(n111), .B(n586), .O(n585));
  orx  g0524(.A(n587), .B(n1109), .O(n586));
  andx g0525(.A(n588), .B(n1124), .O(n587));
  andx g0526(.A(n590), .B(n589), .O(n588));
  invx g0527(.A(n896), .O(n589));
  orx  g0528(.A(n1113), .B(n591), .O(n590));
  orx  g0529(.A(n1226), .B(n592), .O(n591));
  andx g0530(.A(n593), .B(n1242), .O(n592));
  orx  g0531(.A(n594), .B(n82), .O(n593));
  andx g0532(.A(n93), .B(n595), .O(n594));
  orx  g0533(.A(n596), .B(n65), .O(n595));
  andx g0534(.A(n134), .B(n597), .O(n596));
  orx  g0535(.A(n128), .B(n598), .O(n597));
  andx g0536(.A(pi01), .B(n1261), .O(n598));
  invx g0537(.A(n69), .O(n599));
  andx g0538(.A(n601), .B(n150), .O(po19));
  orx  g0539(.A(n602), .B(n1173), .O(n601));
  andx g0540(.A(n1313), .B(n603), .O(n602));
  orx  g0541(.A(n1317), .B(n604), .O(n603));
  andx g0542(.A(n759), .B(n605), .O(n604));
  orx  g0543(.A(n606), .B(n70), .O(n605));
  andx g0544(.A(n648), .B(n607), .O(n606));
  orx  g0545(.A(n608), .B(n1194), .O(n607));
  andx g0546(.A(n1084), .B(n609), .O(n608));
  orx  g0547(.A(n610), .B(n108), .O(n609));
  andx g0548(.A(n611), .B(n1203), .O(n610));
  orx  g0549(.A(n612), .B(n91), .O(n611));
  andx g0550(.A(n960), .B(n613), .O(n612));
  orx  g0551(.A(n616), .B(n614), .O(n613));
  orx  g0552(.A(n72), .B(n615), .O(n614));
  andx g0553(.A(n1032), .B(n99), .O(n615));
  andx g0554(.A(n1032), .B(n617), .O(n616));
  orx  g0555(.A(n618), .B(n80), .O(n617));
  andx g0556(.A(n1028), .B(n619), .O(n618));
  orx  g0557(.A(n1018), .B(n620), .O(n619));
  orx  g0558(.A(n1233), .B(n621), .O(n620));
  andx g0559(.A(n622), .B(n125), .O(n621));
  orx  g0560(.A(n625), .B(n623), .O(n622));
  orx  g0561(.A(n624), .B(n1238), .O(n623));
  andx g0562(.A(n1122), .B(n142), .O(n624));
  andx g0563(.A(n1121), .B(n626), .O(n625));
  orx  g0564(.A(n1252), .B(n627), .O(n626));
  orx  g0565(.A(n629), .B(n628), .O(n627));
  andx g0566(.A(n1250), .B(n1267), .O(n628));
  andx g0567(.A(n1265), .B(n630), .O(n629));
  orx  g0568(.A(n631), .B(n64), .O(n630));
  andx g0569(.A(n109), .B(pi19), .O(n631));
  andx g0570(.A(n633), .B(n153), .O(po18));
  orx  g0571(.A(n634), .B(n1164), .O(n633));
  andx g0572(.A(n724), .B(n635), .O(n634));
  orx  g0573(.A(n1140), .B(n636), .O(n635));
  orx  g0574(.A(n100), .B(n637), .O(n636));
  andx g0575(.A(n1313), .B(n638), .O(n637));
  orx  g0576(.A(n639), .B(n86), .O(n638));
  andx g0577(.A(n640), .B(n131), .O(n639));
  orx  g0578(.A(n641), .B(n1135), .O(n640));
  andx g0579(.A(n759), .B(n642), .O(n641));
  orx  g0580(.A(n643), .B(n1002), .O(n642));
  andx g0581(.A(n1310), .B(n644), .O(n643));
  orx  g0582(.A(n647), .B(n645), .O(n644));
  orx  g0583(.A(n646), .B(n1132), .O(n645));
  andx g0584(.A(n648), .B(n1318), .O(n646));
  andx g0585(.A(n649), .B(n648), .O(n647));
  invx g0586(.A(n1195), .O(n648));
  andx g0587(.A(n650), .B(n1085), .O(n649));
  orx  g0588(.A(n1304), .B(n651), .O(n650));
  andx g0589(.A(n1129), .B(n652), .O(n651));
  orx  g0590(.A(n124), .B(n653), .O(n652));
  andx g0591(.A(n654), .B(n1203), .O(n653));
  orx  g0592(.A(n655), .B(n1094), .O(n654));
  andx g0593(.A(n960), .B(n656), .O(n655));
  orx  g0594(.A(n657), .B(n101), .O(n656));
  andx g0595(.A(n658), .B(n699), .O(n657));
  orx  g0596(.A(n659), .B(n1283), .O(n658));
  andx g0597(.A(n1032), .B(n660), .O(n659));
  orx  g0598(.A(n663), .B(n661), .O(n660));
  orx  g0599(.A(n662), .B(n947), .O(n661));
  andx g0600(.A(n905), .B(n1030), .O(n662));
  andx g0601(.A(n1028), .B(n664), .O(n663));
  orx  g0602(.A(n129), .B(n665), .O(n664));
  andx g0603(.A(n666), .B(n1225), .O(n665));
  orx  g0604(.A(n667), .B(n68), .O(n666));
  andx g0605(.A(n1121), .B(n668), .O(n667));
  orx  g0606(.A(n65), .B(n669), .O(n668));
  andx g0607(.A(n109), .B(pi18), .O(n669));
  andx g0608(.A(n671), .B(n152), .O(po17));
  orx  g0609(.A(n672), .B(n107), .O(n671));
  andx g0610(.A(n1065), .B(n673), .O(n672));
  orx  g0611(.A(n674), .B(n1170), .O(n673));
  andx g0612(.A(n724), .B(n675), .O(n674));
  orx  g0613(.A(n676), .B(n1140), .O(n675));
  andx g0614(.A(n677), .B(n1185), .O(n676));
  orx  g0615(.A(n678), .B(n116), .O(n677));
  andx g0616(.A(n1313), .B(n679), .O(n678));
  orx  g0617(.A(n680), .B(n103), .O(n679));
  andx g0618(.A(n681), .B(n131), .O(n680));
  orx  g0619(.A(n682), .B(n1132), .O(n681));
  andx g0620(.A(n1130), .B(n683), .O(n682));
  orx  g0621(.A(n684), .B(n71), .O(n683));
  andx g0622(.A(n685), .B(n1085), .O(n684));
  orx  g0623(.A(n686), .B(n967), .O(n685));
  andx g0624(.A(n687), .B(n96), .O(n686));
  orx  g0625(.A(n690), .B(n688), .O(n687));
  orx  g0626(.A(n689), .B(n883), .O(n688));
  andx g0627(.A(n964), .B(n123), .O(n689));
  andx g0628(.A(n691), .B(n1203), .O(n690));
  orx  g0629(.A(n692), .B(n67), .O(n691));
  andx g0630(.A(n1292), .B(n693), .O(n692));
  orx  g0631(.A(n696), .B(n694), .O(n693));
  orx  g0632(.A(n695), .B(n831), .O(n694));
  andx g0633(.A(n1096), .B(n149), .O(n695));
  andx g0634(.A(n960), .B(n697), .O(n696));
  orx  g0635(.A(n698), .B(n1103), .O(n697));
  andx g0636(.A(n700), .B(n699), .O(n698));
  invx g0637(.A(n1286), .O(n699));
  orx  g0638(.A(n701), .B(n906), .O(n700));
  andx g0639(.A(n1282), .B(n702), .O(n701));
  orx  g0640(.A(n705), .B(n703), .O(n702));
  orx  g0641(.A(n704), .B(n99), .O(n703));
  andx g0642(.A(n905), .B(n112), .O(n704));
  andx g0643(.A(n1124), .B(n706), .O(n705));
  orx  g0644(.A(n707), .B(n130), .O(n706));
  andx g0645(.A(n708), .B(n1232), .O(n707));
  orx  g0646(.A(n709), .B(n68), .O(n708));
  andx g0647(.A(n1122), .B(n710), .O(n709));
  orx  g0648(.A(n711), .B(n1244), .O(n710));
  andx g0649(.A(n712), .B(n73), .O(n711));
  orx  g0650(.A(n1262), .B(pi17), .O(n712));
  andx g0651(.A(n714), .B(n151), .O(po16));
  orx  g0652(.A(n715), .B(n92), .O(n714));
  andx g0653(.A(n1333), .B(n716), .O(n715));
  orx  g0654(.A(n717), .B(n75), .O(n716));
  andx g0655(.A(n1065), .B(n718), .O(n717));
  orx  g0656(.A(n719), .B(n138), .O(n718));
  andx g0657(.A(n1038), .B(n720), .O(n719));
  orx  g0658(.A(n723), .B(n721), .O(n720));
  orx  g0659(.A(n722), .B(n137), .O(n721));
  andx g0660(.A(n724), .B(pi30), .O(n722));
  andx g0661(.A(n725), .B(n724), .O(n723));
  invx g0662(.A(n1173), .O(n724));
  andx g0663(.A(n726), .B(n1185), .O(n725));
  orx  g0664(.A(n1315), .B(n727), .O(n726));
  andx g0665(.A(n1137), .B(n728), .O(n727));
  orx  g0666(.A(n133), .B(n729), .O(n728));
  andx g0667(.A(n759), .B(n730), .O(n729));
  orx  g0668(.A(n731), .B(n70), .O(n730));
  andx g0669(.A(n1131), .B(n732), .O(n731));
  orx  g0670(.A(n733), .B(n110), .O(n732));
  andx g0671(.A(n734), .B(n801), .O(n733));
  andx g0672(.A(n758), .B(n735), .O(n734));
  orx  g0673(.A(n736), .B(n67), .O(n735));
  andx g0674(.A(n1287), .B(n737), .O(n736));
  orx  g0675(.A(n738), .B(n961), .O(n737));
  andx g0676(.A(n1101), .B(n739), .O(n738));
  orx  g0677(.A(n740), .B(n906), .O(n739));
  andx g0678(.A(n1032), .B(n741), .O(n740));
  orx  g0679(.A(n742), .B(n99), .O(n741));
  andx g0680(.A(n851), .B(n743), .O(n742));
  orx  g0681(.A(n744), .B(n80), .O(n743));
  andx g0682(.A(n1029), .B(n745), .O(n744));
  orx  g0683(.A(n746), .B(n1219), .O(n745));
  andx g0684(.A(n747), .B(n1228), .O(n746));
  andx g0685(.A(n748), .B(n125), .O(n747));
  orx  g0686(.A(n749), .B(n68), .O(n748));
  andx g0687(.A(n959), .B(n750), .O(n749));
  orx  g0688(.A(n751), .B(n105), .O(n750));
  andx g0689(.A(n752), .B(n1242), .O(n751));
  orx  g0690(.A(n753), .B(n1245), .O(n752));
  andx g0691(.A(n81), .B(n754), .O(n753));
  orx  g0692(.A(n755), .B(n847), .O(n754));
  andx g0693(.A(n904), .B(n756), .O(n755));
  orx  g0694(.A(pi16), .B(n757), .O(n756));
  invx g0695(.A(n1260), .O(n757));
  invx g0696(.A(n74), .O(n758));
  invx g0697(.A(n1077), .O(n759));
  andx g0698(.A(n761), .B(n150), .O(po15));
  orx  g0699(.A(n762), .B(n1147), .O(n761));
  andx g0700(.A(n908), .B(n763), .O(n762));
  orx  g0701(.A(n764), .B(n1339), .O(n763));
  andx g0702(.A(n1333), .B(n765), .O(n764));
  orx  g0703(.A(n766), .B(n1160), .O(n765));
  andx g0704(.A(n852), .B(n767), .O(n766));
  orx  g0705(.A(n768), .B(n1063), .O(n767));
  andx g0706(.A(n1325), .B(n769), .O(n768));
  orx  g0707(.A(n770), .B(n120), .O(n769));
  andx g0708(.A(n1181), .B(n771), .O(n770));
  orx  g0709(.A(n772), .B(n100), .O(n771));
  andx g0710(.A(n803), .B(n773), .O(n772));
  orx  g0711(.A(n774), .B(n140), .O(n773));
  andx g0712(.A(n1137), .B(n775), .O(n774));
  orx  g0713(.A(n776), .B(n103), .O(n775));
  andx g0714(.A(n1134), .B(n777), .O(n776));
  orx  g0715(.A(n778), .B(n98), .O(n777));
  andx g0716(.A(n1310), .B(n779), .O(n778));
  orx  g0717(.A(n780), .B(n110), .O(n779));
  andx g0718(.A(n801), .B(n781), .O(n780));
  orx  g0719(.A(n782), .B(n74), .O(n781));
  andx g0720(.A(n1128), .B(n783), .O(n782));
  orx  g0721(.A(n784), .B(n831), .O(n783));
  andx g0722(.A(n1287), .B(n785), .O(n784));
  orx  g0723(.A(n786), .B(n148), .O(n785));
  andx g0724(.A(n960), .B(n787), .O(n786));
  orx  g0725(.A(n791), .B(n788), .O(n787));
  orx  g0726(.A(n789), .B(n1099), .O(n788));
  andx g0727(.A(n790), .B(n1283), .O(n789));
  invx g0728(.A(n906), .O(n790));
  andx g0729(.A(n1127), .B(n792), .O(n791));
  orx  g0730(.A(n793), .B(n892), .O(n792));
  andx g0731(.A(n794), .B(n1228), .O(n793));
  andx g0732(.A(n795), .B(n1225), .O(n794));
  orx  g0733(.A(n1233), .B(n796), .O(n795));
  andx g0734(.A(n1270), .B(n797), .O(n796));
  orx  g0735(.A(n798), .B(n94), .O(n797));
  andx g0736(.A(n1265), .B(n799), .O(n798));
  orx  g0737(.A(n800), .B(n64), .O(n799));
  andx g0738(.A(pi15), .B(n109), .O(n800));
  invx g0739(.A(n802), .O(n801));
  orx  g0740(.A(n79), .B(n71), .O(n802));
  invx g0741(.A(n116), .O(n803));
  andx g0742(.A(n805), .B(n153), .O(po14));
  orx  g0743(.A(n806), .B(n1358), .O(n805));
  andx g0744(.A(n1146), .B(n807), .O(n806));
  orx  g0745(.A(n78), .B(n808), .O(n807));
  orx  g0746(.A(n810), .B(n809), .O(n808));
  andx g0747(.A(n908), .B(n145), .O(n809));
  andx g0748(.A(n1338), .B(n811), .O(n810));
  orx  g0749(.A(n812), .B(n102), .O(n811));
  andx g0750(.A(n1333), .B(n813), .O(n812));
  orx  g0751(.A(n814), .B(n117), .O(n813));
  andx g0752(.A(n852), .B(n815), .O(n814));
  orx  g0753(.A(n816), .B(n138), .O(n815));
  andx g0754(.A(n1175), .B(n817), .O(n816));
  orx  g0755(.A(pi30), .B(n818), .O(n817));
  andx g0756(.A(n819), .B(n1182), .O(n818));
  orx  g0757(.A(n1315), .B(n820), .O(n819));
  andx g0758(.A(n1134), .B(n821), .O(n820));
  orx  g0759(.A(n822), .B(n1194), .O(n821));
  andx g0760(.A(n1300), .B(n823), .O(n822));
  orx  g0761(.A(n824), .B(n79), .O(n823));
  andx g0762(.A(n966), .B(n825), .O(n824));
  orx  g0763(.A(n826), .B(n74), .O(n825));
  andx g0764(.A(n1128), .B(n827), .O(n826));
  orx  g0765(.A(n833), .B(n828), .O(n827));
  orx  g0766(.A(n829), .B(n1293), .O(n828));
  andx g0767(.A(n830), .B(n91), .O(n829));
  invx g0768(.A(n831), .O(n830));
  orx  g0769(.A(n832), .B(n1293), .O(n831));
  andx g0770(.A(n1355), .B(n148), .O(n832));
  andx g0771(.A(n1287), .B(n834), .O(n833));
  orx  g0772(.A(n835), .B(n1283), .O(n834));
  andx g0773(.A(n1032), .B(n836), .O(n835));
  orx  g0774(.A(n837), .B(n99), .O(n836));
  andx g0775(.A(n851), .B(n838), .O(n837));
  orx  g0776(.A(n839), .B(n112), .O(n838));
  andx g0777(.A(n136), .B(n840), .O(n839));
  orx  g0778(.A(n841), .B(n1125), .O(n840));
  andx g0779(.A(n842), .B(n66), .O(n841));
  orx  g0780(.A(n843), .B(n896), .O(n842));
  andx g0781(.A(n844), .B(n125), .O(n843));
  orx  g0782(.A(n845), .B(n68), .O(n844));
  andx g0783(.A(n959), .B(n846), .O(n845));
  orx  g0784(.A(n849), .B(n847), .O(n846));
  orx  g0785(.A(n848), .B(n63), .O(n847));
  andx g0786(.A(n93), .B(n65), .O(n848));
  andx g0787(.A(n850), .B(n73), .O(n849));
  orx  g0788(.A(n1262), .B(pi14), .O(n850));
  invx g0789(.A(n947), .O(n851));
  invx g0790(.A(n75), .O(n852));
  andx g0791(.A(n854), .B(n1357), .O(po13));
  andx g0792(.A(n1040), .B(n855), .O(n854));
  orx  g0793(.A(n856), .B(n1045), .O(n855));
  andx g0794(.A(n1146), .B(n857), .O(n856));
  orx  g0795(.A(n858), .B(n90), .O(n857));
  andx g0796(.A(n1349), .B(n859), .O(n858));
  orx  g0797(.A(n860), .B(n1053), .O(n859));
  andx g0798(.A(n908), .B(n861), .O(n860));
  orx  g0799(.A(n862), .B(n119), .O(n861));
  andx g0800(.A(n863), .B(n144), .O(n862));
  orx  g0801(.A(n864), .B(n1343), .O(n863));
  andx g0802(.A(n1141), .B(n865), .O(n864));
  orx  g0803(.A(n867), .B(n75), .O(n865));
  orx  g0804(.A(n1341), .B(n117), .O(n866));
  andx g0805(.A(n1325), .B(n868), .O(n867));
  orx  g0806(.A(n871), .B(n869), .O(n868));
  orx  g0807(.A(n870), .B(n120), .O(n869));
  andx g0808(.A(n1038), .B(n137), .O(n870));
  andx g0809(.A(n872), .B(n1365), .O(n871));
  orx  g0810(.A(n140), .B(n873), .O(n872));
  andx g0811(.A(n1137), .B(n874), .O(n873));
  orx  g0812(.A(n875), .B(n103), .O(n874));
  andx g0813(.A(n876), .B(n131), .O(n875));
  orx  g0814(.A(n877), .B(n1002), .O(n876));
  andx g0815(.A(n1130), .B(n878), .O(n877));
  orx  g0816(.A(n879), .B(n83), .O(n878));
  andx g0817(.A(n880), .B(n1301), .O(n879));
  orx  g0818(.A(n881), .B(n967), .O(n880));
  andx g0819(.A(n882), .B(n96), .O(n881));
  orx  g0820(.A(n885), .B(n883), .O(n882));
  orx  g0821(.A(n884), .B(n74), .O(n883));
  andx g0822(.A(n1129), .B(n1296), .O(n884));
  andx g0823(.A(n1129), .B(n886), .O(n885));
  orx  g0824(.A(n887), .B(n964), .O(n886));
  andx g0825(.A(n1292), .B(n888), .O(n887));
  orx  g0826(.A(n889), .B(n906), .O(n888));
  orx  g0827(.A(n890), .B(n91), .O(n889));
  andx g0828(.A(n905), .B(n891), .O(n890));
  orx  g0829(.A(n894), .B(n892), .O(n891));
  orx  g0830(.A(n893), .B(n1278), .O(n892));
  andx g0831(.A(n136), .B(n1307), .O(n893));
  andx g0832(.A(n136), .B(n895), .O(n894));
  orx  g0833(.A(n897), .B(n896), .O(n895));
  andx g0834(.A(n1226), .B(pi19), .O(n896));
  andx g0835(.A(n898), .B(n125), .O(n897));
  orx  g0836(.A(n899), .B(n1238), .O(n898));
  andx g0837(.A(n1122), .B(n900), .O(n899));
  orx  g0838(.A(n901), .B(n82), .O(n900));
  andx g0839(.A(n904), .B(n902), .O(n901));
  orx  g0840(.A(n903), .B(n127), .O(n902));
  andx g0841(.A(pi13), .B(n1261), .O(n903));
  invx g0842(.A(n64), .O(n904));
  invx g0843(.A(n80), .O(n905));
  orx  g0844(.A(n72), .B(n907), .O(n906));
  andx g0845(.A(n1106), .B(pi19), .O(n907));
  invx g0846(.A(n92), .O(n908));
  orx  g0847(.A(n911), .B(n910), .O(po12));
  andx g0848(.A(n1042), .B(n152), .O(n910));
  andx g0849(.A(n1356), .B(n912), .O(n911));
  orx  g0850(.A(n913), .B(n1353), .O(n912));
  andx g0851(.A(n1044), .B(n914), .O(n913));
  orx  g0852(.A(n917), .B(n915), .O(n914));
  orx  g0853(.A(n916), .B(n1045), .O(n915));
  andx g0854(.A(pi18), .B(n1362), .O(n916));
  andx g0855(.A(n89), .B(n918), .O(n917));
  orx  g0856(.A(n919), .B(n76), .O(n918));
  andx g0857(.A(n969), .B(n920), .O(n919));
  orx  g0858(.A(n119), .B(n921), .O(n920));
  orx  g0859(.A(n1337), .B(n922), .O(n921));
  andx g0860(.A(n1141), .B(n923), .O(n922));
  orx  g0861(.A(n924), .B(n117), .O(n923));
  andx g0862(.A(n87), .B(n925), .O(n924));
  orx  g0863(.A(n928), .B(n926), .O(n925));
  orx  g0864(.A(n927), .B(n120), .O(n926));
  andx g0865(.A(n1038), .B(pi30), .O(n927));
  andx g0866(.A(n1038), .B(n929), .O(n928));
  orx  g0867(.A(n930), .B(n1183), .O(n929));
  andx g0868(.A(n931), .B(n1185), .O(n930));
  orx  g0869(.A(n932), .B(n116), .O(n931));
  andx g0870(.A(n1137), .B(n933), .O(n932));
  orx  g0871(.A(n934), .B(n997), .O(n933));
  andx g0872(.A(n935), .B(n1001), .O(n934));
  andx g0873(.A(n966), .B(n936), .O(n935));
  orx  g0874(.A(n937), .B(n108), .O(n936));
  andx g0875(.A(n1295), .B(n938), .O(n937));
  orx  g0876(.A(n939), .B(n124), .O(n938));
  andx g0877(.A(n963), .B(n940), .O(n939));
  orx  g0878(.A(n84), .B(n941), .O(n940));
  andx g0879(.A(n1128), .B(n942), .O(n941));
  orx  g0880(.A(n943), .B(n1094), .O(n942));
  andx g0881(.A(n960), .B(n944), .O(n943));
  orx  g0882(.A(n1286), .B(n945), .O(n944));
  andx g0883(.A(n1282), .B(n946), .O(n945));
  orx  g0884(.A(n949), .B(n947), .O(n946));
  orx  g0885(.A(n948), .B(n1279), .O(n947));
  andx g0886(.A(n1166), .B(n130), .O(n948));
  andx g0887(.A(n1029), .B(n950), .O(n949));
  orx  g0888(.A(n951), .B(n112), .O(n950));
  andx g0889(.A(n136), .B(n952), .O(n951));
  orx  g0890(.A(n1223), .B(n953), .O(n952));
  orx  g0891(.A(n1233), .B(n954), .O(n953));
  andx g0892(.A(n959), .B(n955), .O(n954));
  orx  g0893(.A(n956), .B(n1244), .O(n955));
  andx g0894(.A(n1265), .B(n957), .O(n956));
  orx  g0895(.A(n958), .B(n64), .O(n957));
  andx g0896(.A(pi12), .B(n1260), .O(n958));
  invx g0897(.A(n1238), .O(n959));
  invx g0898(.A(n961), .O(n960));
  orx  g0899(.A(n962), .B(n148), .O(n961));
  andx g0900(.A(n1106), .B(n113), .O(n962));
  invx g0901(.A(n964), .O(n963));
  orx  g0902(.A(n965), .B(n124), .O(n964));
  andx g0903(.A(n1166), .B(n149), .O(n965));
  invx g0904(.A(n967), .O(n966));
  orx  g0905(.A(n968), .B(n79), .O(n967));
  andx g0906(.A(pi18), .B(n97), .O(n968));
  invx g0907(.A(n1053), .O(n969));
  andx g0908(.A(n1040), .B(n971), .O(po11));
  orx  g0909(.A(n972), .B(n1359), .O(n971));
  andx g0910(.A(n1357), .B(n973), .O(n972));
  orx  g0911(.A(n974), .B(n104), .O(n973));
  andx g0912(.A(n1352), .B(n975), .O(n974));
  orx  g0913(.A(n982), .B(n976), .O(n975));
  orx  g0914(.A(n1049), .B(n977), .O(n976));
  orx  g0915(.A(n981), .B(n978), .O(n977));
  andx g0916(.A(n1146), .B(n76), .O(n978));
  orx  g0917(.A(n980), .B(n1153), .O(n979));
  andx g0918(.A(n1330), .B(n146), .O(n980));
  andx g0919(.A(n1349), .B(n1053), .O(n981));
  andx g0920(.A(n1143), .B(n983), .O(n982));
  orx  g0921(.A(n985), .B(n984), .O(n983));
  orx  g0922(.A(n1363), .B(n1337), .O(n984));
  andx g0923(.A(n1039), .B(n986), .O(n985));
  orx  g0924(.A(n989), .B(n987), .O(n986));
  orx  g0925(.A(n988), .B(n107), .O(n987));
  andx g0926(.A(n1285), .B(pi30), .O(n988));
  andx g0927(.A(n87), .B(n990), .O(n989));
  orx  g0928(.A(n991), .B(n69), .O(n990));
  andx g0929(.A(n1038), .B(n992), .O(n991));
  orx  g0930(.A(n993), .B(n137), .O(n992));
  andx g0931(.A(n1181), .B(n994), .O(n993));
  orx  g0932(.A(n995), .B(n1071), .O(n994));
  andx g0933(.A(n1035), .B(n996), .O(n995));
  orx  g0934(.A(n1000), .B(n997), .O(n996));
  orx  g0935(.A(n998), .B(n1077), .O(n997));
  andx g0936(.A(n1001), .B(n71), .O(n998));
  orx  g0937(.A(n83), .B(n1302), .O(n999));
  andx g0938(.A(n1004), .B(n1001), .O(n1000));
  invx g0939(.A(n1002), .O(n1001));
  orx  g0940(.A(n1003), .B(n1077), .O(n1002));
  andx g0941(.A(n1285), .B(n1318), .O(n1003));
  andx g0942(.A(n1005), .B(n96), .O(n1004));
  orx  g0943(.A(n1006), .B(n1296), .O(n1005));
  andx g0944(.A(n1007), .B(n123), .O(n1006));
  orx  g0945(.A(n1206), .B(n1008), .O(n1007));
  andx g0946(.A(n1128), .B(n1009), .O(n1008));
  orx  g0947(.A(n1306), .B(n1010), .O(n1009));
  andx g0948(.A(n1034), .B(n1011), .O(n1010));
  orx  g0949(.A(n1012), .B(n101), .O(n1011));
  andx g0950(.A(n1032), .B(n1013), .O(n1012));
  orx  g0951(.A(n1014), .B(n99), .O(n1013));
  andx g0952(.A(n1029), .B(n1015), .O(n1014));
  orx  g0953(.A(n1016), .B(n112), .O(n1015));
  andx g0954(.A(n1028), .B(n1017), .O(n1016));
  orx  g0955(.A(n1019), .B(n1018), .O(n1017));
  orx  g0956(.A(n1110), .B(n95), .O(n1018));
  andx g0957(.A(n1123), .B(n1020), .O(n1019));
  orx  g0958(.A(n126), .B(n1021), .O(n1020));
  andx g0959(.A(n1270), .B(n1022), .O(n1021));
  orx  g0960(.A(n1023), .B(n105), .O(n1022));
  andx g0961(.A(n1024), .B(n1242), .O(n1023));
  orx  g0962(.A(n65), .B(n1025), .O(n1024));
  andx g0963(.A(n1265), .B(n1026), .O(n1025));
  orx  g0964(.A(n1027), .B(n64), .O(n1026));
  andx g0965(.A(pi11), .B(n1260), .O(n1027));
  invx g0966(.A(n1220), .O(n1028));
  invx g0967(.A(n1030), .O(n1029));
  orx  g0968(.A(n1031), .B(n80), .O(n1030));
  andx g0969(.A(n1330), .B(n129), .O(n1031));
  invx g0970(.A(n85), .O(n1032));
  orx  g0971(.A(n1106), .B(n1283), .O(n1033));
  invx g0972(.A(n1103), .O(n1034));
  invx g0973(.A(n103), .O(n1035));
  orx  g0974(.A(n1037), .B(n86), .O(n1036));
  andx g0975(.A(pi19), .B(n132), .O(n1037));
  invx g0976(.A(n1170), .O(n1038));
  invx g0977(.A(n102), .O(n1039));
  andx g0978(.A(n153), .B(n1041), .O(n1040));
  invx g0979(.A(n1042), .O(n1041));
  andx g0980(.A(n1359), .B(pi18), .O(n1042));
  andx g0981(.A(n1047), .B(n1044), .O(po10));
  invx g0982(.A(n1045), .O(n1044));
  orx  g0983(.A(n1046), .B(n104), .O(n1045));
  andx g0984(.A(pi19), .B(n1362), .O(n1046));
  andx g0985(.A(n1048), .B(n151), .O(n1047));
  orx  g0986(.A(n1051), .B(n1049), .O(n1048));
  orx  g0987(.A(n1050), .B(n122), .O(n1049));
  andx g0988(.A(n1146), .B(n1153), .O(n1050));
  andx g0989(.A(n1146), .B(n1052), .O(n1051));
  orx  g0990(.A(n1055), .B(n1053), .O(n1052));
  orx  g0991(.A(n1054), .B(n78), .O(n1053));
  andx g0992(.A(n1355), .B(n146), .O(n1054));
  andx g0993(.A(n1143), .B(n1056), .O(n1055));
  orx  g0994(.A(n1057), .B(n1339), .O(n1056));
  andx g0995(.A(n1142), .B(n1058), .O(n1057));
  orx  g0996(.A(n1061), .B(n102), .O(n1058));
  orx  g0997(.A(n1060), .B(n1343), .O(n1059));
  andx g0998(.A(n1341), .B(pi20), .O(n1060));
  andx g0999(.A(n1141), .B(n1062), .O(n1061));
  orx  g1000(.A(n1066), .B(n1063), .O(n1062));
  orx  g1001(.A(n1064), .B(n1331), .O(n1063));
  andx g1002(.A(n1065), .B(n69), .O(n1064));
  invx g1003(.A(n1164), .O(n1065));
  andx g1004(.A(n1325), .B(n1067), .O(n1066));
  orx  g1005(.A(n1068), .B(n1169), .O(n1067));
  andx g1006(.A(n1175), .B(n1069), .O(n1068));
  orx  g1007(.A(n1140), .B(n1070), .O(n1069));
  orx  g1008(.A(n1073), .B(n1071), .O(n1070));
  orx  g1009(.A(n1072), .B(n116), .O(n1071));
  andx g1010(.A(n1314), .B(n139), .O(n1072));
  andx g1011(.A(n1137), .B(n1074), .O(n1073));
  orx  g1012(.A(n1317), .B(n1075), .O(n1074));
  andx g1013(.A(n1134), .B(n1076), .O(n1075));
  orx  g1014(.A(n1079), .B(n1077), .O(n1076));
  orx  g1015(.A(n1078), .B(n133), .O(n1077));
  andx g1016(.A(n1336), .B(n83), .O(n1078));
  andx g1017(.A(n1131), .B(n1080), .O(n1079));
  orx  g1018(.A(n1086), .B(n1081), .O(n1080));
  orx  g1019(.A(n1082), .B(n1195), .O(n1081));
  andx g1020(.A(n1130), .B(n1083), .O(n1082));
  invx g1021(.A(n1084), .O(n1083));
  andx g1022(.A(n1085), .B(n1319), .O(n1084));
  invx g1023(.A(n79), .O(n1085));
  andx g1024(.A(n1130), .B(n1087), .O(n1086));
  orx  g1025(.A(n1090), .B(n74), .O(n1087));
  orx  g1026(.A(n1089), .B(n97), .O(n1088));
  andx g1027(.A(n1305), .B(n1355), .O(n1089));
  andx g1028(.A(n1129), .B(n1091), .O(n1090));
  orx  g1029(.A(n84), .B(n1092), .O(n1091));
  andx g1030(.A(n1128), .B(n1093), .O(n1092));
  orx  g1031(.A(n1097), .B(n1094), .O(n1093));
  orx  g1032(.A(n1095), .B(n1293), .O(n1094));
  andx g1033(.A(n1096), .B(n118), .O(n1095));
  invx g1034(.A(n91), .O(n1096));
  andx g1035(.A(n1098), .B(n147), .O(n1097));
  orx  g1036(.A(n1107), .B(n1099), .O(n1098));
  orx  g1037(.A(n1100), .B(n1103), .O(n1099));
  andx g1038(.A(n1101), .B(n72), .O(n1100));
  invx g1039(.A(n101), .O(n1101));
  orx  g1040(.A(n1105), .B(n1103), .O(n1102));
  orx  g1041(.A(n1104), .B(n149), .O(n1103));
  andx g1042(.A(n1345), .B(n1307), .O(n1104));
  andx g1043(.A(n1106), .B(pi20), .O(n1105));
  andx g1044(.A(n129), .B(n1342), .O(n1106));
  andx g1045(.A(n1127), .B(n1108), .O(n1107));
  orx  g1046(.A(n1111), .B(n1109), .O(n1108));
  orx  g1047(.A(n1110), .B(n1220), .O(n1109));
  andx g1048(.A(n130), .B(n1124), .O(n1110));
  andx g1049(.A(n1123), .B(n1112), .O(n1111));
  orx  g1050(.A(n1114), .B(n1113), .O(n1112));
  andx g1051(.A(n68), .B(n125), .O(n1113));
  andx g1052(.A(n1122), .B(n1115), .O(n1114));
  orx  g1053(.A(n1116), .B(n143), .O(n1115));
  andx g1054(.A(n1121), .B(n1117), .O(n1116));
  orx  g1055(.A(n1118), .B(n94), .O(n1117));
  andx g1056(.A(n1265), .B(n1119), .O(n1118));
  orx  g1057(.A(n127), .B(n1120), .O(n1119));
  andx g1058(.A(pi10), .B(n1261), .O(n1120));
  invx g1059(.A(n1245), .O(n1121));
  invx g1060(.A(n105), .O(n1122));
  andx g1061(.A(n1225), .B(n1124), .O(n1123));
  invx g1062(.A(n1125), .O(n1124));
  orx  g1063(.A(n1126), .B(n95), .O(n1125));
  andx g1064(.A(pi18), .B(n130), .O(n1126));
  invx g1065(.A(n1279), .O(n1127));
  invx g1066(.A(n67), .O(n1128));
  invx g1067(.A(n108), .O(n1129));
  invx g1068(.A(n1194), .O(n1130));
  invx g1069(.A(n1132), .O(n1131));
  orx  g1070(.A(n1133), .B(n70), .O(n1132));
  andx g1071(.A(n114), .B(n83), .O(n1133));
  invx g1072(.A(n1135), .O(n1134));
  orx  g1073(.A(n1136), .B(n132), .O(n1135));
  andx g1074(.A(n1345), .B(n1318), .O(n1136));
  invx g1075(.A(n86), .O(n1137));
  orx  g1076(.A(n1139), .B(n140), .O(n1138));
  andx g1077(.A(pi20), .B(n132), .O(n1139));
  invx g1078(.A(n1181), .O(n1140));
  invx g1079(.A(n1160), .O(n1141));
  invx g1080(.A(n1343), .O(n1142));
  invx g1081(.A(n119), .O(n1143));
  orx  g1082(.A(n1145), .B(n92), .O(n1144));
  andx g1083(.A(pi18), .B(n145), .O(n1145));
  invx g1084(.A(n1147), .O(n1146));
  orx  g1085(.A(n1148), .B(n122), .O(n1147));
  andx g1086(.A(n1166), .B(n145), .O(n1148));
  andx g1087(.A(n1356), .B(n1150), .O(po00));
  orx  g1088(.A(n1151), .B(n104), .O(n1150));
  andx g1089(.A(n1352), .B(n1152), .O(n1151));
  orx  g1090(.A(n1155), .B(n90), .O(n1152));
  orx  g1091(.A(n1154), .B(n122), .O(n1153));
  andx g1092(.A(n113), .B(n146), .O(n1154));
  andx g1093(.A(n1349), .B(n1156), .O(n1155));
  orx  g1094(.A(n92), .B(n1157), .O(n1156));
  orx  g1095(.A(n1337), .B(n1158), .O(n1157));
  andx g1096(.A(n1333), .B(n1159), .O(n1158));
  orx  g1097(.A(n1162), .B(n1160), .O(n1159));
  orx  g1098(.A(n1161), .B(n107), .O(n1160));
  andx g1099(.A(n1341), .B(pi19), .O(n1161));
  andx g1100(.A(n87), .B(n1163), .O(n1162));
  orx  g1101(.A(n1167), .B(n1164), .O(n1163));
  orx  g1102(.A(n1165), .B(n88), .O(n1164));
  andx g1103(.A(n1166), .B(pi30), .O(n1165));
  andx g1104(.A(pi18), .B(n114), .O(n1166));
  andx g1105(.A(n1325), .B(n1168), .O(n1167));
  orx  g1106(.A(n1180), .B(n1169), .O(n1168));
  orx  g1107(.A(n1172), .B(n1170), .O(n1169));
  orx  g1108(.A(n1171), .B(n120), .O(n1170));
  andx g1109(.A(n1355), .B(pi30), .O(n1171));
  andx g1110(.A(n1175), .B(n1173), .O(n1172));
  orx  g1111(.A(n1174), .B(n137), .O(n1173));
  andx g1112(.A(pi18), .B(pi30), .O(n1174));
  invx g1113(.A(n137), .O(n1175));
  orx  g1114(.A(n1179), .B(n120), .O(n1176));
  orx  g1115(.A(n1178), .B(n1331), .O(n1177));
  andx g1116(.A(pi30), .B(pi20), .O(n1178));
  andx g1117(.A(pi19), .B(pi30), .O(n1179));
  andx g1118(.A(n1184), .B(n1181), .O(n1180));
  andx g1119(.A(n1182), .B(n1365), .O(n1181));
  invx g1120(.A(n1183), .O(n1182));
  andx g1121(.A(n100), .B(pi19), .O(n1183));
  andx g1122(.A(n1186), .B(n1185), .O(n1184));
  invx g1123(.A(n100), .O(n1185));
  orx  g1124(.A(n1190), .B(n116), .O(n1186));
  orx  g1125(.A(n1189), .B(n100), .O(n1187));
  andx g1126(.A(n140), .B(pi20), .O(n1188));
  andx g1127(.A(pi19), .B(n140), .O(n1189));
  andx g1128(.A(n1313), .B(n1191), .O(n1190));
  orx  g1129(.A(n1317), .B(n1192), .O(n1191));
  andx g1130(.A(n1310), .B(n1193), .O(n1192));
  orx  g1131(.A(n1198), .B(n1194), .O(n1193));
  orx  g1132(.A(n1197), .B(n1195), .O(n1194));
  orx  g1133(.A(n1196), .B(n70), .O(n1195));
  andx g1134(.A(pi20), .B(n83), .O(n1196));
  andx g1135(.A(pi19), .B(n1318), .O(n1197));
  andx g1136(.A(n1300), .B(n1199), .O(n1198));
  orx  g1137(.A(n1200), .B(n108), .O(n1199));
  andx g1138(.A(n1295), .B(n1201), .O(n1200));
  orx  g1139(.A(n1202), .B(n1305), .O(n1201));
  andx g1140(.A(n1204), .B(n1203), .O(n1202));
  invx g1141(.A(n1206), .O(n1203));
  orx  g1142(.A(n1209), .B(n67), .O(n1204));
  orx  g1143(.A(n1208), .B(n1206), .O(n1205));
  orx  g1144(.A(n1207), .B(n124), .O(n1206));
  andx g1145(.A(n114), .B(n148), .O(n1207));
  andx g1146(.A(n1330), .B(n148), .O(n1208));
  andx g1147(.A(n1292), .B(n1210), .O(n1209));
  orx  g1148(.A(n1211), .B(n91), .O(n1210));
  andx g1149(.A(n1287), .B(n1212), .O(n1211));
  orx  g1150(.A(n1286), .B(n1213), .O(n1212));
  andx g1151(.A(n1282), .B(n1214), .O(n1213));
  orx  g1152(.A(n1217), .B(n80), .O(n1214));
  orx  g1153(.A(n1216), .B(n1279), .O(n1215));
  andx g1154(.A(n113), .B(n129), .O(n1216));
  andx g1155(.A(n111), .B(n1218), .O(n1217));
  orx  g1156(.A(n1227), .B(n1219), .O(n1218));
  orx  g1157(.A(n1222), .B(n1220), .O(n1219));
  orx  g1158(.A(n1221), .B(n1278), .O(n1220));
  andx g1159(.A(n1355), .B(n1307), .O(n1221));
  andx g1160(.A(n1228), .B(n1223), .O(n1222));
  invx g1161(.A(n1224), .O(n1223));
  andx g1162(.A(n66), .B(n1225), .O(n1224));
  invx g1163(.A(n1226), .O(n1225));
  andx g1164(.A(n126), .B(pi20), .O(n1226));
  andx g1165(.A(n1231), .B(n1228), .O(n1227));
  invx g1166(.A(n95), .O(n1228));
  orx  g1167(.A(n1230), .B(n112), .O(n1229));
  andx g1168(.A(pi19), .B(n130), .O(n1230));
  andx g1169(.A(n1234), .B(n1232), .O(n1231));
  invx g1170(.A(n1233), .O(n1232));
  andx g1171(.A(n1272), .B(pi19), .O(n1233));
  orx  g1172(.A(n1235), .B(n1272), .O(n1234));
  andx g1173(.A(n1270), .B(n1236), .O(n1235));
  orx  g1174(.A(n1241), .B(n105), .O(n1236));
  orx  g1175(.A(n1240), .B(n1238), .O(n1237));
  orx  g1176(.A(n1239), .B(n126), .O(n1238));
  andx g1177(.A(n143), .B(pi20), .O(n1239));
  andx g1178(.A(n1274), .B(pi19), .O(n1240));
  andx g1179(.A(n1243), .B(n1242), .O(n1241));
  invx g1180(.A(n142), .O(n1242));
  orx  g1181(.A(n1255), .B(n1244), .O(n1243));
  orx  g1182(.A(n1247), .B(n1245), .O(n1244));
  orx  g1183(.A(n1246), .B(n143), .O(n1245));
  andx g1184(.A(n1345), .B(n127), .O(n1246));
  andx g1185(.A(n1250), .B(n65), .O(n1247));
  orx  g1186(.A(n1249), .B(n1267), .O(n1248));
  andx g1187(.A(n114), .B(n128), .O(n1249));
  invx g1188(.A(n63), .O(n1250));
  orx  g1189(.A(n1254), .B(n1252), .O(n1251));
  orx  g1190(.A(n1253), .B(n143), .O(n1252));
  andx g1191(.A(n1336), .B(n127), .O(n1253));
  andx g1192(.A(n1285), .B(n128), .O(n1254));
  andx g1193(.A(n1265), .B(n1256), .O(n1255));
  orx  g1194(.A(n1259), .B(n64), .O(n1256));
  orx  g1195(.A(n1258), .B(n1266), .O(n1257));
  andx g1196(.A(pi19), .B(n127), .O(n1258));
  andx g1197(.A(pi00), .B(n1260), .O(n1259));
  andx g1198(.A(n1261), .B(n73), .O(n1260));
  invx g1199(.A(n1262), .O(n1261));
  andx g1200(.A(n1264), .B(n1263), .O(n1262));
  andx g1201(.A(n62), .B(n1336), .O(n1263));
  invx g1202(.A(n1321), .O(n1264));
  invx g1203(.A(n1266), .O(n1265));
  orx  g1204(.A(n1269), .B(n1267), .O(n1266));
  orx  g1205(.A(n1268), .B(n142), .O(n1267));
  andx g1206(.A(pi21), .B(n128), .O(n1268));
  andx g1207(.A(pi20), .B(n127), .O(n1269));
  invx g1208(.A(n68), .O(n1270));
  orx  g1209(.A(n1273), .B(n1272), .O(n1271));
  andx g1210(.A(pi21), .B(n143), .O(n1272));
  andx g1211(.A(n1274), .B(n113), .O(n1273));
  andx g1212(.A(n128), .B(n62), .O(n1274));
  invx g1213(.A(n73), .O(n1275));
  orx  g1214(.A(n1375), .B(n1277), .O(n1276));
  orx  g1215(.A(pi24), .B(n1321), .O(n1277));
  orx  g1216(.A(n1281), .B(n99), .O(n1278));
  orx  g1217(.A(n1280), .B(n1306), .O(n1279));
  andx g1218(.A(pi21), .B(n129), .O(n1280));
  andx g1219(.A(pi20), .B(n1307), .O(n1281));
  invx g1220(.A(n1283), .O(n1282));
  orx  g1221(.A(n1286), .B(n1284), .O(n1283));
  andx g1222(.A(n1285), .B(n130), .O(n1284));
  andx g1223(.A(pi21), .B(pi19), .O(n1285));
  andx g1224(.A(n130), .B(n1336), .O(n1286));
  invx g1225(.A(n118), .O(n1287));
  orx  g1226(.A(n1291), .B(n91), .O(n1288));
  orx  g1227(.A(n1290), .B(n1293), .O(n1289));
  andx g1228(.A(pi19), .B(n149), .O(n1290));
  andx g1229(.A(pi18), .B(n1306), .O(n1291));
  invx g1230(.A(n1293), .O(n1292));
  orx  g1231(.A(n1294), .B(n124), .O(n1293));
  andx g1232(.A(pi20), .B(n1306), .O(n1294));
  invx g1233(.A(n1296), .O(n1295));
  orx  g1234(.A(n1299), .B(n108), .O(n1296));
  orx  g1235(.A(n1298), .B(n97), .O(n1297));
  andx g1236(.A(n124), .B(pi19), .O(n1298));
  andx g1237(.A(n1305), .B(pi18), .O(n1299));
  andx g1238(.A(n1301), .B(n1319), .O(n1300));
  invx g1239(.A(n1302), .O(n1301));
  andx g1240(.A(n79), .B(pi18), .O(n1302));
  andx g1241(.A(n97), .B(pi19), .O(n1303));
  andx g1242(.A(pi20), .B(n1305), .O(n1304));
  andx g1243(.A(n148), .B(pi21), .O(n1305));
  andx g1244(.A(n129), .B(n62), .O(n1306));
  invx g1245(.A(n66), .O(n1307));
  orx  g1246(.A(n1378), .B(n1309), .O(n1308));
  orx  g1247(.A(pi23), .B(n1321), .O(n1309));
  invx g1248(.A(n70), .O(n1310));
  orx  g1249(.A(n1312), .B(n133), .O(n1311));
  andx g1250(.A(pi21), .B(n1318), .O(n1312));
  invx g1251(.A(n1314), .O(n1313));
  orx  g1252(.A(n1316), .B(n1315), .O(n1314));
  andx g1253(.A(n133), .B(pi21), .O(n1315));
  andx g1254(.A(n113), .B(n133), .O(n1316));
  andx g1255(.A(n83), .B(n62), .O(n1317));
  invx g1256(.A(n1319), .O(n1318));
  orx  g1257(.A(n1378), .B(n1320), .O(n1319));
  orx  g1258(.A(n1321), .B(n1375), .O(n1320));
  orx  g1259(.A(n1323), .B(n1322), .O(n1321));
  orx  g1260(.A(n1370), .B(n1369), .O(n1322));
  orx  g1261(.A(n1372), .B(n1324), .O(n1323));
  orx  g1262(.A(n1377), .B(n1373), .O(n1324));
  invx g1263(.A(n138), .O(n1325));
  orx  g1264(.A(n1329), .B(n69), .O(n1326));
  orx  g1265(.A(n1328), .B(n1331), .O(n1327));
  andx g1266(.A(n114), .B(pi30), .O(n1328));
  andx g1267(.A(n1330), .B(pi30), .O(n1329));
  andx g1268(.A(pi20), .B(pi18), .O(n1330));
  orx  g1269(.A(n1332), .B(n145), .O(n1331));
  andx g1270(.A(pi21), .B(pi30), .O(n1332));
  invx g1271(.A(n107), .O(n1333));
  orx  g1272(.A(n1335), .B(n146), .O(n1334));
  andx g1273(.A(n1336), .B(pi30), .O(n1335));
  andx g1274(.A(pi20), .B(pi21), .O(n1336));
  andx g1275(.A(n1343), .B(n1338), .O(n1337));
  invx g1276(.A(n1339), .O(n1338));
  orx  g1277(.A(n1340), .B(n1363), .O(n1339));
  andx g1278(.A(n1341), .B(n114), .O(n1340));
  andx g1279(.A(pi30), .B(n1342), .O(n1341));
  andx g1280(.A(pi21), .B(pi18), .O(n1342));
  orx  g1281(.A(n1344), .B(n145), .O(n1343));
  andx g1282(.A(n1345), .B(pi30), .O(n1344));
  andx g1283(.A(pi21), .B(n113), .O(n1345));
  andx g1284(.A(pi20), .B(pi19), .O(n1346));
  orx  g1285(.A(n1348), .B(n78), .O(n1347));
  andx g1286(.A(pi19), .B(n1363), .O(n1348));
  invx g1287(.A(n78), .O(n1349));
  orx  g1288(.A(n1351), .B(n122), .O(n1350));
  andx g1289(.A(pi20), .B(n1363), .O(n1351));
  invx g1290(.A(n1353), .O(n1352));
  orx  g1291(.A(n1354), .B(n104), .O(n1353));
  andx g1292(.A(n1355), .B(n122), .O(n1354));
  andx g1293(.A(pi19), .B(pi18), .O(n1355));
  andx g1294(.A(n152), .B(n1357), .O(n1356));
  invx g1295(.A(n1358), .O(n1357));
  orx  g1296(.A(n1360), .B(n1359), .O(n1358));
  andx g1297(.A(n1361), .B(pi19), .O(n1359));
  andx g1298(.A(pi18), .B(n1361), .O(n1360));
  andx g1299(.A(pi20), .B(n1362), .O(n1361));
  andx g1300(.A(n146), .B(pi21), .O(n1362));
  andx g1301(.A(n62), .B(pi30), .O(n1363));
  orx  g1302(.A(n1366), .B(n1365), .O(n1364));
  invx g1303(.A(pi30), .O(n1365));
  andx g1304(.A(n1374), .B(n1367), .O(n1366));
  andx g1305(.A(n1371), .B(n1368), .O(n1367));
  andx g1306(.A(n1370), .B(n1369), .O(n1368));
  invx g1307(.A(pi29), .O(n1369));
  invx g1308(.A(pi28), .O(n1370));
  andx g1309(.A(n1373), .B(n1372), .O(n1371));
  invx g1310(.A(pi27), .O(n1372));
  invx g1311(.A(pi26), .O(n1373));
  andx g1312(.A(n1376), .B(n1375), .O(n1374));
  invx g1313(.A(pi23), .O(n1375));
  andx g1314(.A(n1378), .B(n1377), .O(n1376));
  invx g1315(.A(pi25), .O(n1377));
  invx g1316(.A(pi24), .O(n1378));
endmodule


