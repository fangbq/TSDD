// Benchmark "top" written by ABC on Fri Feb  7 13:34:28 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21;
  wire n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n874, n875, n876, n877, n878, n879, n880, n882, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1023, n1024, n1026, n1027,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1274, n1275,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
    n1328;
  invx g0000(.a(pi40), .O(n72));
  andx g0001(.a(pi44), .b(n72), .O(n73));
  invx g0002(.a(pi43), .O(n74));
  andx g0003(.a(n74), .b(pi45), .O(n75));
  andx g0004(.a(n75), .b(n73), .O(n76));
  andx g0005(.a(n76), .b(pi46), .O(n77));
  andx g0006(.a(pi43), .b(pi44), .O(n78));
  invx g0007(.a(pi44), .O(n79));
  andx g0008(.a(pi43), .b(n79), .O(n80));
  andx g0009(.a(n80), .b(pi40), .O(n81));
  andx g0010(.a(n81), .b(pi37), .O(n82));
  orx  g0011(.a(n82), .b(n78), .O(n83));
  andx g0012(.a(n74), .b(pi40), .O(n84));
  orx  g0013(.a(n84), .b(n83), .O(n85));
  invx g0014(.a(n85), .O(n86));
  andx g0015(.a(n86), .b(pi22), .O(n87));
  invx g0016(.a(pi22), .O(n88));
  andx g0017(.a(pi44), .b(pi40), .O(n89));
  andx g0018(.a(n89), .b(n74), .O(n90));
  andx g0019(.a(n90), .b(n88), .O(n91));
  andx g0020(.a(n88), .b(pi40), .O(n92));
  invx g0021(.a(n92), .O(n93));
  andx g0022(.a(pi19), .b(pi37), .O(n94));
  invx g0023(.a(pi37), .O(n95));
  andx g0024(.a(pi28), .b(n95), .O(n96));
  orx  g0025(.a(n96), .b(pi40), .O(n97));
  orx  g0026(.a(n97), .b(n94), .O(n98));
  andx g0027(.a(n98), .b(n93), .O(n99));
  andx g0028(.a(n99), .b(n83), .O(n100));
  orx  g0029(.a(n100), .b(n91), .O(n101));
  orx  g0030(.a(n101), .b(n87), .O(n102));
  invx g0031(.a(n102), .O(n103));
  invx g0032(.a(pi32), .O(n104));
  orx  g0033(.a(n74), .b(n79), .O(n105));
  andx g0034(.a(pi37), .b(pi27), .O(n106));
  orx  g0035(.a(n106), .b(n105), .O(n107));
  andx g0036(.a(pi39), .b(n95), .O(n108));
  andx g0037(.a(n108), .b(pi25), .O(n109));
  invx g0038(.a(n109), .O(n110));
  andx g0039(.a(pi16), .b(pi37), .O(n111));
  invx g0040(.a(n111), .O(n112));
  invx g0041(.a(pi29), .O(n113));
  orx  g0042(.a(pi39), .b(pi37), .O(n114));
  orx  g0043(.a(n114), .b(n113), .O(n115));
  andx g0044(.a(n115), .b(n112), .O(n116));
  andx g0045(.a(n116), .b(n110), .O(n117));
  orx  g0046(.a(n117), .b(n107), .O(n118));
  orx  g0047(.a(pi24), .b(pi27), .O(n119));
  andx g0048(.a(n119), .b(n74), .O(n120));
  invx g0049(.a(n120), .O(n121));
  andx g0050(.a(n121), .b(n107), .O(n122));
  andx g0051(.a(n122), .b(pi21), .O(n123));
  andx g0052(.a(n107), .b(pi23), .O(n124));
  andx g0053(.a(n124), .b(n120), .O(n125));
  orx  g0054(.a(n125), .b(n123), .O(n126));
  invx g0055(.a(n126), .O(n127));
  andx g0056(.a(n127), .b(n118), .O(n128));
  invx g0057(.a(n128), .O(n129));
  andx g0058(.a(n129), .b(n104), .O(n130));
  invx g0059(.a(pi35), .O(n131));
  andx g0060(.a(n128), .b(n131), .O(n132));
  orx  g0061(.a(n132), .b(n130), .O(n133));
  orx  g0062(.a(n133), .b(n103), .O(n134));
  orx  g0063(.a(n134), .b(n77), .O(n135));
  invx g0064(.a(pi16), .O(n136));
  invx g0065(.a(n89), .O(n137));
  andx g0066(.a(n137), .b(n95), .O(n138));
  orx  g0067(.a(n138), .b(pi43), .O(n139));
  invx g0068(.a(n139), .O(n140));
  orx  g0069(.a(n140), .b(n83), .O(n141));
  orx  g0070(.a(n141), .b(n136), .O(n142));
  andx g0071(.a(pi16), .b(pi40), .O(n143));
  andx g0072(.a(n90), .b(n136), .O(n144));
  invx g0073(.a(n144), .O(n145));
  orx  g0074(.a(n74), .b(pi44), .O(n146));
  orx  g0075(.a(n146), .b(n72), .O(n147));
  orx  g0076(.a(n147), .b(n95), .O(n148));
  andx g0077(.a(n148), .b(n105), .O(n149));
  andx g0078(.a(pi15), .b(pi37), .O(n150));
  invx g0079(.a(n150), .O(n151));
  invx g0080(.a(pi19), .O(n152));
  orx  g0081(.a(n152), .b(pi37), .O(n153));
  andx g0082(.a(n153), .b(n72), .O(n154));
  andx g0083(.a(n154), .b(n151), .O(n155));
  orx  g0084(.a(n155), .b(n149), .O(n156));
  andx g0085(.a(n156), .b(n145), .O(n157));
  orx  g0086(.a(n157), .b(n143), .O(n158));
  andx g0087(.a(n158), .b(n142), .O(n159));
  invx g0088(.a(pi20), .O(n160));
  orx  g0089(.a(n114), .b(n160), .O(n161));
  invx g0090(.a(pi17), .O(n162));
  invx g0091(.a(pi39), .O(n163));
  orx  g0092(.a(n163), .b(pi37), .O(n164));
  orx  g0093(.a(n164), .b(n162), .O(n165));
  andx g0094(.a(pi10), .b(pi37), .O(n166));
  invx g0095(.a(n166), .O(n167));
  andx g0096(.a(n167), .b(n165), .O(n168));
  andx g0097(.a(n168), .b(n161), .O(n169));
  orx  g0098(.a(n169), .b(n107), .O(n170));
  invx g0099(.a(pi23), .O(n171));
  invx g0100(.a(pi27), .O(n172));
  orx  g0101(.a(n95), .b(n172), .O(n173));
  andx g0102(.a(n173), .b(n78), .O(n174));
  orx  g0103(.a(n174), .b(n171), .O(n175));
  invx g0104(.a(pi24), .O(n176));
  orx  g0105(.a(n176), .b(pi43), .O(n177));
  orx  g0106(.a(n177), .b(pi27), .O(n178));
  orx  g0107(.a(n178), .b(n175), .O(n179));
  invx g0108(.a(pi11), .O(n180));
  andx g0109(.a(pi24), .b(n74), .O(n181));
  andx g0110(.a(n181), .b(n172), .O(n182));
  orx  g0111(.a(n182), .b(n174), .O(n183));
  orx  g0112(.a(n183), .b(n180), .O(n184));
  andx g0113(.a(n184), .b(n179), .O(n185));
  andx g0114(.a(n185), .b(n170), .O(n186));
  orx  g0115(.a(n186), .b(n104), .O(n187));
  invx g0116(.a(n161), .O(n188));
  andx g0117(.a(n108), .b(pi17), .O(n189));
  orx  g0118(.a(n166), .b(n189), .O(n190));
  orx  g0119(.a(n190), .b(n188), .O(n191));
  andx g0120(.a(n191), .b(n174), .O(n192));
  andx g0121(.a(n182), .b(n124), .O(n193));
  andx g0122(.a(n178), .b(n107), .O(n194));
  andx g0123(.a(n194), .b(pi11), .O(n195));
  orx  g0124(.a(n195), .b(n193), .O(n196));
  orx  g0125(.a(n196), .b(n192), .O(n197));
  orx  g0126(.a(n197), .b(n131), .O(n198));
  andx g0127(.a(n198), .b(n187), .O(n199));
  orx  g0128(.a(n199), .b(n159), .O(n200));
  orx  g0129(.a(n114), .b(n162), .O(n201));
  invx g0130(.a(n201), .O(n202));
  andx g0131(.a(n108), .b(pi11), .O(n203));
  andx g0132(.a(pi06), .b(pi37), .O(n204));
  orx  g0133(.a(n204), .b(n203), .O(n205));
  orx  g0134(.a(n205), .b(n202), .O(n206));
  andx g0135(.a(n206), .b(n174), .O(n207));
  andx g0136(.a(n194), .b(pi12), .O(n208));
  orx  g0137(.a(n208), .b(n193), .O(n209));
  orx  g0138(.a(n209), .b(n207), .O(n210));
  orx  g0139(.a(n210), .b(n131), .O(n211));
  orx  g0140(.a(n164), .b(n180), .O(n212));
  invx g0141(.a(n204), .O(n213));
  andx g0142(.a(n213), .b(n212), .O(n214));
  andx g0143(.a(n214), .b(n201), .O(n215));
  orx  g0144(.a(n215), .b(n107), .O(n216));
  invx g0145(.a(pi12), .O(n217));
  orx  g0146(.a(n183), .b(n217), .O(n218));
  andx g0147(.a(n218), .b(n179), .O(n219));
  andx g0148(.a(n219), .b(n216), .O(n220));
  orx  g0149(.a(n220), .b(n104), .O(n221));
  andx g0150(.a(n221), .b(n211), .O(n222));
  invx g0151(.a(pi15), .O(n223));
  orx  g0152(.a(n141), .b(n223), .O(n224));
  andx g0153(.a(n90), .b(n223), .O(n225));
  invx g0154(.a(n225), .O(n226));
  andx g0155(.a(n223), .b(pi40), .O(n227));
  andx g0156(.a(pi13), .b(pi37), .O(n228));
  invx g0157(.a(n228), .O(n229));
  invx g0158(.a(pi18), .O(n230));
  orx  g0159(.a(n230), .b(pi37), .O(n231));
  andx g0160(.a(n231), .b(n72), .O(n232));
  andx g0161(.a(n232), .b(n229), .O(n233));
  orx  g0162(.a(n233), .b(n227), .O(n234));
  orx  g0163(.a(n234), .b(n149), .O(n235));
  andx g0164(.a(n235), .b(n226), .O(n236));
  andx g0165(.a(n236), .b(n224), .O(n237));
  orx  g0166(.a(n237), .b(n222), .O(n238));
  invx g0167(.a(pi31), .O(n239));
  andx g0168(.a(n186), .b(n239), .O(n240));
  invx g0169(.a(pi30), .O(n241));
  andx g0170(.a(n197), .b(n241), .O(n242));
  orx  g0171(.a(n242), .b(n240), .O(n243));
  andx g0172(.a(n243), .b(n159), .O(n244));
  orx  g0173(.a(n244), .b(n238), .O(n245));
  andx g0174(.a(n245), .b(n200), .O(n246));
  andx g0175(.a(n108), .b(pi20), .O(n247));
  invx g0176(.a(n114), .O(n248));
  andx g0177(.a(n248), .b(pi21), .O(n249));
  orx  g0178(.a(n249), .b(n228), .O(n250));
  orx  g0179(.a(n250), .b(n247), .O(n251));
  andx g0180(.a(n251), .b(n174), .O(n252));
  andx g0181(.a(n194), .b(pi17), .O(n253));
  orx  g0182(.a(n253), .b(n193), .O(n254));
  orx  g0183(.a(n254), .b(n252), .O(n255));
  invx g0184(.a(n255), .O(n256));
  andx g0185(.a(n256), .b(pi31), .O(n257));
  andx g0186(.a(n139), .b(n149), .O(n258));
  andx g0187(.a(n258), .b(pi18), .O(n259));
  andx g0188(.a(n90), .b(n230), .O(n260));
  andx g0189(.a(pi22), .b(n95), .O(n261));
  orx  g0190(.a(n261), .b(pi40), .O(n262));
  orx  g0191(.a(n262), .b(n111), .O(n263));
  andx g0192(.a(n136), .b(n230), .O(n264));
  andx g0193(.a(pi16), .b(pi18), .O(n265));
  orx  g0194(.a(n265), .b(n264), .O(n266));
  orx  g0195(.a(n266), .b(n72), .O(n267));
  andx g0196(.a(n267), .b(n263), .O(n268));
  andx g0197(.a(n268), .b(n83), .O(n269));
  orx  g0198(.a(n269), .b(n260), .O(n270));
  orx  g0199(.a(n270), .b(n259), .O(n271));
  andx g0200(.a(n255), .b(pi30), .O(n272));
  orx  g0201(.a(n272), .b(n271), .O(n273));
  orx  g0202(.a(n273), .b(n257), .O(n274));
  invx g0203(.a(n274), .O(n275));
  orx  g0204(.a(n275), .b(n246), .O(n276));
  invx g0205(.a(n271), .O(n277));
  andx g0206(.a(n255), .b(n104), .O(n278));
  orx  g0207(.a(n255), .b(pi35), .O(n279));
  invx g0208(.a(n279), .O(n280));
  orx  g0209(.a(n280), .b(n278), .O(n281));
  orx  g0210(.a(n281), .b(n277), .O(n282));
  andx g0211(.a(n282), .b(n276), .O(n283));
  andx g0212(.a(n108), .b(pi21), .O(n284));
  andx g0213(.a(n248), .b(pi25), .O(n285));
  orx  g0214(.a(n285), .b(n150), .O(n286));
  orx  g0215(.a(n286), .b(n284), .O(n287));
  andx g0216(.a(n287), .b(n174), .O(n288));
  andx g0217(.a(n177), .b(n160), .O(n289));
  andx g0218(.a(n181), .b(n171), .O(n290));
  orx  g0219(.a(n290), .b(n289), .O(n291));
  orx  g0220(.a(n291), .b(n174), .O(n292));
  invx g0221(.a(n292), .O(n293));
  orx  g0222(.a(n293), .b(n288), .O(n294));
  invx g0223(.a(n294), .O(n295));
  andx g0224(.a(n295), .b(pi31), .O(n296));
  invx g0225(.a(n296), .O(n297));
  andx g0226(.a(n258), .b(pi19), .O(n298));
  invx g0227(.a(n298), .O(n299));
  andx g0228(.a(n90), .b(n152), .O(n300));
  invx g0229(.a(n300), .O(n301));
  andx g0230(.a(n264), .b(n152), .O(n302));
  andx g0231(.a(n302), .b(pi40), .O(n303));
  invx g0232(.a(pi26), .O(n304));
  andx g0233(.a(pi37), .b(n72), .O(n305));
  orx  g0234(.a(n305), .b(n304), .O(n306));
  andx g0235(.a(pi18), .b(pi37), .O(n307));
  orx  g0236(.a(n307), .b(pi40), .O(n308));
  invx g0237(.a(n308), .O(n309));
  andx g0238(.a(n309), .b(n306), .O(n310));
  orx  g0239(.a(n310), .b(n303), .O(n311));
  orx  g0240(.a(n311), .b(n149), .O(n312));
  andx g0241(.a(n312), .b(n301), .O(n313));
  andx g0242(.a(n313), .b(n299), .O(n314));
  andx g0243(.a(n294), .b(pi30), .O(n315));
  invx g0244(.a(n315), .O(n316));
  andx g0245(.a(n316), .b(n314), .O(n317));
  andx g0246(.a(n317), .b(n297), .O(n318));
  orx  g0247(.a(n318), .b(n283), .O(n319));
  andx g0248(.a(n294), .b(n104), .O(n320));
  orx  g0249(.a(n294), .b(pi35), .O(n321));
  invx g0250(.a(n321), .O(n322));
  orx  g0251(.a(n322), .b(n320), .O(n323));
  orx  g0252(.a(n323), .b(n314), .O(n324));
  andx g0253(.a(n324), .b(n319), .O(n325));
  orx  g0254(.a(n325), .b(n77), .O(n326));
  invx g0255(.a(n134), .O(n327));
  andx g0256(.a(n102), .b(n77), .O(n328));
  invx g0257(.a(n328), .O(n329));
  andx g0258(.a(n128), .b(pi31), .O(n330));
  andx g0259(.a(n129), .b(pi30), .O(n331));
  orx  g0260(.a(n331), .b(n102), .O(n332));
  orx  g0261(.a(n332), .b(n330), .O(n333));
  andx g0262(.a(n333), .b(n329), .O(n334));
  orx  g0263(.a(n334), .b(n327), .O(n335));
  andx g0264(.a(n335), .b(n135), .O(n336));
  invx g0265(.a(n336), .O(n337));
  orx  g0266(.a(n337), .b(n326), .O(n338));
  andx g0267(.a(n338), .b(n135), .O(n339));
  andx g0268(.a(n258), .b(pi15), .O(n340));
  invx g0269(.a(n227), .O(n341));
  andx g0270(.a(pi18), .b(n95), .O(n342));
  orx  g0271(.a(n342), .b(pi40), .O(n343));
  orx  g0272(.a(n343), .b(n228), .O(n344));
  andx g0273(.a(n344), .b(n341), .O(n345));
  andx g0274(.a(n345), .b(n83), .O(n346));
  orx  g0275(.a(n346), .b(n225), .O(n347));
  orx  g0276(.a(n347), .b(n340), .O(n348));
  andx g0277(.a(n210), .b(pi30), .O(n349));
  andx g0278(.a(n220), .b(pi31), .O(n350));
  orx  g0279(.a(n350), .b(n349), .O(n351));
  orx  g0280(.a(n351), .b(n348), .O(n352));
  andx g0281(.a(n352), .b(n238), .O(n353));
  andx g0282(.a(n258), .b(pi16), .O(n354));
  invx g0283(.a(n143), .O(n355));
  andx g0284(.a(pi19), .b(n95), .O(n356));
  orx  g0285(.a(n356), .b(pi40), .O(n357));
  orx  g0286(.a(n357), .b(n150), .O(n358));
  andx g0287(.a(n358), .b(n83), .O(n359));
  orx  g0288(.a(n359), .b(n144), .O(n360));
  andx g0289(.a(n360), .b(n355), .O(n361));
  orx  g0290(.a(n361), .b(n354), .O(n362));
  orx  g0291(.a(n197), .b(pi31), .O(n363));
  orx  g0292(.a(n186), .b(pi30), .O(n364));
  andx g0293(.a(n364), .b(n363), .O(n365));
  orx  g0294(.a(n365), .b(n362), .O(n366));
  andx g0295(.a(n366), .b(n200), .O(n367));
  andx g0296(.a(n367), .b(n353), .O(n368));
  invx g0297(.a(n313), .O(n369));
  orx  g0298(.a(n369), .b(n298), .O(n370));
  orx  g0299(.a(n315), .b(n370), .O(n371));
  orx  g0300(.a(n371), .b(n296), .O(n372));
  andx g0301(.a(n324), .b(n372), .O(n373));
  andx g0302(.a(n282), .b(n274), .O(n374));
  andx g0303(.a(n374), .b(n373), .O(n375));
  andx g0304(.a(n375), .b(n368), .O(n376));
  orx  g0305(.a(n376), .b(n77), .O(n377));
  andx g0306(.a(n220), .b(pi35), .O(n378));
  andx g0307(.a(n295), .b(n256), .O(n379));
  andx g0308(.a(n379), .b(n186), .O(n380));
  andx g0309(.a(n380), .b(n378), .O(n381));
  invx g0310(.a(n77), .O(n382));
  andx g0311(.a(n210), .b(n131), .O(n383));
  andx g0312(.a(n255), .b(n197), .O(n384));
  andx g0313(.a(n384), .b(n294), .O(n385));
  andx g0314(.a(n385), .b(n383), .O(n386));
  orx  g0315(.a(n386), .b(n382), .O(n387));
  orx  g0316(.a(n387), .b(n381), .O(n388));
  andx g0317(.a(n388), .b(pi14), .O(n389));
  andx g0318(.a(n389), .b(n377), .O(n390));
  andx g0319(.a(n390), .b(n336), .O(n391));
  andx g0320(.a(n86), .b(pi26), .O(n392));
  invx g0321(.a(n392), .O(n393));
  andx g0322(.a(pi22), .b(pi37), .O(n394));
  andx g0323(.a(pi33), .b(n95), .O(n395));
  orx  g0324(.a(n395), .b(n394), .O(n396));
  andx g0325(.a(n396), .b(n72), .O(n397));
  andx g0326(.a(n397), .b(n83), .O(n398));
  invx g0327(.a(n398), .O(n399));
  andx g0328(.a(n137), .b(n148), .O(n400));
  orx  g0329(.a(n400), .b(pi26), .O(n401));
  andx g0330(.a(n401), .b(n399), .O(n402));
  andx g0331(.a(n402), .b(n393), .O(n403));
  invx g0332(.a(n403), .O(n404));
  andx g0333(.a(n404), .b(n77), .O(n405));
  invx g0334(.a(n405), .O(n406));
  andx g0335(.a(n108), .b(pi29), .O(n407));
  andx g0336(.a(n248), .b(pi34), .O(n408));
  orx  g0337(.a(n408), .b(n307), .O(n409));
  orx  g0338(.a(n409), .b(n407), .O(n410));
  andx g0339(.a(n410), .b(n174), .O(n411));
  andx g0340(.a(n122), .b(pi25), .O(n412));
  orx  g0341(.a(n412), .b(n125), .O(n413));
  orx  g0342(.a(n413), .b(n411), .O(n414));
  andx g0343(.a(n414), .b(n104), .O(n415));
  invx g0344(.a(n415), .O(n416));
  orx  g0345(.a(n414), .b(pi35), .O(n417));
  andx g0346(.a(n417), .b(n416), .O(n418));
  andx g0347(.a(n418), .b(n404), .O(n419));
  invx g0348(.a(n419), .O(n420));
  invx g0349(.a(n414), .O(n421));
  andx g0350(.a(n421), .b(pi31), .O(n422));
  andx g0351(.a(n414), .b(pi30), .O(n423));
  orx  g0352(.a(n423), .b(n404), .O(n424));
  orx  g0353(.a(n424), .b(n422), .O(n425));
  andx g0354(.a(n425), .b(n420), .O(n426));
  andx g0355(.a(n426), .b(n406), .O(n427));
  andx g0356(.a(n419), .b(n77), .O(n428));
  orx  g0357(.a(n428), .b(n427), .O(n429));
  orx  g0358(.a(n429), .b(n391), .O(n430));
  invx g0359(.a(n368), .O(n431));
  invx g0360(.a(n320), .O(n432));
  andx g0361(.a(n321), .b(n432), .O(n433));
  andx g0362(.a(n433), .b(n370), .O(n434));
  orx  g0363(.a(n434), .b(n318), .O(n435));
  invx g0364(.a(n278), .O(n436));
  andx g0365(.a(n279), .b(n436), .O(n437));
  andx g0366(.a(n437), .b(n271), .O(n438));
  orx  g0367(.a(n438), .b(n275), .O(n439));
  orx  g0368(.a(n439), .b(n435), .O(n440));
  orx  g0369(.a(n440), .b(n431), .O(n441));
  andx g0370(.a(n441), .b(n382), .O(n442));
  invx g0371(.a(n389), .O(n443));
  orx  g0372(.a(n443), .b(n442), .O(n444));
  orx  g0373(.a(n444), .b(n337), .O(n445));
  invx g0374(.a(n429), .O(n446));
  orx  g0375(.a(n446), .b(n445), .O(n447));
  andx g0376(.a(n447), .b(n430), .O(n448));
  andx g0377(.a(n448), .b(n339), .O(n449));
  invx g0378(.a(n135), .O(n450));
  andx g0379(.a(n197), .b(pi32), .O(n451));
  andx g0380(.a(n186), .b(pi35), .O(n452));
  orx  g0381(.a(n452), .b(n451), .O(n453));
  andx g0382(.a(n453), .b(n362), .O(n454));
  andx g0383(.a(n210), .b(pi32), .O(n455));
  orx  g0384(.a(n455), .b(n378), .O(n456));
  andx g0385(.a(n348), .b(n456), .O(n457));
  andx g0386(.a(n366), .b(n457), .O(n458));
  orx  g0387(.a(n458), .b(n454), .O(n459));
  andx g0388(.a(n274), .b(n459), .O(n460));
  orx  g0389(.a(n438), .b(n460), .O(n461));
  andx g0390(.a(n372), .b(n461), .O(n462));
  orx  g0391(.a(n434), .b(n462), .O(n463));
  andx g0392(.a(n463), .b(n382), .O(n464));
  andx g0393(.a(n336), .b(n464), .O(n465));
  orx  g0394(.a(n465), .b(n450), .O(n466));
  andx g0395(.a(n446), .b(n445), .O(n467));
  andx g0396(.a(n429), .b(n391), .O(n468));
  orx  g0397(.a(n468), .b(n467), .O(n469));
  andx g0398(.a(n469), .b(n466), .O(n470));
  orx  g0399(.a(n470), .b(n449), .O(n471));
  orx  g0400(.a(n390), .b(n464), .O(n472));
  andx g0401(.a(n86), .b(pi28), .O(n473));
  invx g0402(.a(pi28), .O(n474));
  andx g0403(.a(n474), .b(n304), .O(n475));
  andx g0404(.a(pi28), .b(pi26), .O(n476));
  orx  g0405(.a(n476), .b(n475), .O(n477));
  andx g0406(.a(n477), .b(pi40), .O(n478));
  andx g0407(.a(n305), .b(pi26), .O(n479));
  andx g0408(.a(n95), .b(n72), .O(n480));
  andx g0409(.a(n480), .b(pi36), .O(n481));
  orx  g0410(.a(n481), .b(n479), .O(n482));
  orx  g0411(.a(n482), .b(n478), .O(n483));
  andx g0412(.a(n483), .b(n83), .O(n484));
  andx g0413(.a(n90), .b(n474), .O(n485));
  orx  g0414(.a(n485), .b(n484), .O(n486));
  orx  g0415(.a(n486), .b(n473), .O(n487));
  invx g0416(.a(n487), .O(n488));
  andx g0417(.a(n108), .b(pi34), .O(n489));
  andx g0418(.a(n248), .b(pi42), .O(n490));
  orx  g0419(.a(n490), .b(n94), .O(n491));
  orx  g0420(.a(n491), .b(n489), .O(n492));
  andx g0421(.a(n492), .b(n174), .O(n493));
  andx g0422(.a(n122), .b(pi29), .O(n494));
  orx  g0423(.a(n494), .b(n125), .O(n495));
  orx  g0424(.a(n495), .b(n493), .O(n496));
  andx g0425(.a(n496), .b(n104), .O(n497));
  invx g0426(.a(n496), .O(n498));
  andx g0427(.a(n498), .b(n131), .O(n499));
  orx  g0428(.a(n499), .b(n497), .O(n500));
  orx  g0429(.a(n500), .b(n488), .O(n501));
  andx g0430(.a(n501), .b(n333), .O(n502));
  andx g0431(.a(n498), .b(pi31), .O(n503));
  andx g0432(.a(n496), .b(pi30), .O(n504));
  orx  g0433(.a(n504), .b(n487), .O(n505));
  orx  g0434(.a(n505), .b(n503), .O(n506));
  andx g0435(.a(n506), .b(n134), .O(n507));
  andx g0436(.a(n507), .b(n502), .O(n508));
  andx g0437(.a(n108), .b(pi42), .O(n509));
  andx g0438(.a(n248), .b(pi48), .O(n510));
  orx  g0439(.a(n510), .b(n394), .O(n511));
  orx  g0440(.a(n511), .b(n509), .O(n512));
  andx g0441(.a(n512), .b(n174), .O(n513));
  andx g0442(.a(n122), .b(pi34), .O(n514));
  orx  g0443(.a(n514), .b(n125), .O(n515));
  orx  g0444(.a(n515), .b(n513), .O(n516));
  invx g0445(.a(n516), .O(n517));
  andx g0446(.a(n517), .b(pi31), .O(n518));
  andx g0447(.a(n86), .b(pi33), .O(n519));
  invx g0448(.a(n519), .O(n520));
  invx g0449(.a(pi33), .O(n521));
  andx g0450(.a(n475), .b(n521), .O(n522));
  orx  g0451(.a(n522), .b(n72), .O(n523));
  andx g0452(.a(n305), .b(pi28), .O(n524));
  andx g0453(.a(n480), .b(pi38), .O(n525));
  orx  g0454(.a(n525), .b(n524), .O(n526));
  invx g0455(.a(n526), .O(n527));
  andx g0456(.a(n527), .b(n523), .O(n528));
  orx  g0457(.a(n528), .b(n149), .O(n529));
  andx g0458(.a(n90), .b(n521), .O(n530));
  invx g0459(.a(n530), .O(n531));
  andx g0460(.a(n531), .b(n529), .O(n532));
  andx g0461(.a(n532), .b(n520), .O(n533));
  invx g0462(.a(n533), .O(n534));
  andx g0463(.a(n516), .b(pi30), .O(n535));
  orx  g0464(.a(n535), .b(n534), .O(n536));
  orx  g0465(.a(n536), .b(n518), .O(n537));
  andx g0466(.a(n516), .b(n104), .O(n538));
  andx g0467(.a(n517), .b(n131), .O(n539));
  orx  g0468(.a(n539), .b(n538), .O(n540));
  orx  g0469(.a(n540), .b(n533), .O(n541));
  andx g0470(.a(n541), .b(n537), .O(n542));
  andx g0471(.a(n542), .b(n426), .O(n543));
  andx g0472(.a(n543), .b(n508), .O(n544));
  andx g0473(.a(n544), .b(n472), .O(n545));
  invx g0474(.a(n541), .O(n546));
  invx g0475(.a(n501), .O(n547));
  andx g0476(.a(n425), .b(n327), .O(n548));
  orx  g0477(.a(n548), .b(n419), .O(n549));
  andx g0478(.a(n549), .b(n506), .O(n550));
  orx  g0479(.a(n550), .b(n547), .O(n551));
  andx g0480(.a(n551), .b(n537), .O(n552));
  orx  g0481(.a(n552), .b(n546), .O(n553));
  orx  g0482(.a(n553), .b(n545), .O(n554));
  invx g0483(.a(n554), .O(n555));
  andx g0484(.a(n555), .b(n471), .O(n556));
  invx g0485(.a(n556), .O(n557));
  andx g0486(.a(n81), .b(n172), .O(n558));
  orx  g0487(.a(n555), .b(n471), .O(n559));
  andx g0488(.a(n559), .b(n558), .O(n560));
  andx g0489(.a(n560), .b(n557), .O(n561));
  andx g0490(.a(n73), .b(pi24), .O(n562));
  orx  g0491(.a(n562), .b(n74), .O(n563));
  andx g0492(.a(n563), .b(n471), .O(n564));
  andx g0493(.a(n95), .b(n79), .O(n565));
  andx g0494(.a(n565), .b(n446), .O(n566));
  invx g0495(.a(n566), .O(n567));
  andx g0496(.a(n104), .b(pi40), .O(n568));
  orx  g0497(.a(n568), .b(n105), .O(n569));
  andx g0498(.a(pi35), .b(pi40), .O(n570));
  andx g0499(.a(n570), .b(pi30), .O(n571));
  andx g0500(.a(n571), .b(pi31), .O(n572));
  andx g0501(.a(n572), .b(pi10), .O(n573));
  andx g0502(.a(n570), .b(n241), .O(n574));
  andx g0503(.a(n574), .b(pi31), .O(n575));
  andx g0504(.a(n575), .b(pi13), .O(n576));
  andx g0505(.a(n239), .b(pi40), .O(n577));
  invx g0506(.a(n570), .O(n578));
  andx g0507(.a(pi30), .b(pi40), .O(n579));
  invx g0508(.a(n579), .O(n580));
  andx g0509(.a(n580), .b(n578), .O(n581));
  andx g0510(.a(n581), .b(n577), .O(n582));
  andx g0511(.a(n582), .b(pi06), .O(n583));
  orx  g0512(.a(n583), .b(n576), .O(n584));
  orx  g0513(.a(n584), .b(n573), .O(n585));
  andx g0514(.a(n571), .b(n239), .O(n586));
  andx g0515(.a(n586), .b(pi15), .O(n587));
  orx  g0516(.a(n587), .b(n95), .O(n588));
  andx g0517(.a(n579), .b(n578), .O(n589));
  andx g0518(.a(n589), .b(pi31), .O(n590));
  andx g0519(.a(n590), .b(pi18), .O(n591));
  invx g0520(.a(n577), .O(n592));
  andx g0521(.a(n581), .b(n592), .O(n593));
  andx g0522(.a(n593), .b(pi19), .O(n594));
  orx  g0523(.a(n594), .b(n591), .O(n595));
  andx g0524(.a(n574), .b(n239), .O(n596));
  andx g0525(.a(n596), .b(pi16), .O(n597));
  andx g0526(.a(n589), .b(n239), .O(n598));
  andx g0527(.a(n598), .b(pi22), .O(n599));
  orx  g0528(.a(n599), .b(n597), .O(n600));
  orx  g0529(.a(n600), .b(n595), .O(n601));
  orx  g0530(.a(n601), .b(n588), .O(n602));
  orx  g0531(.a(n602), .b(n585), .O(n603));
  andx g0532(.a(n586), .b(pi01), .O(n604));
  andx g0533(.a(n572), .b(pi47), .O(n605));
  andx g0534(.a(n575), .b(pi41), .O(n606));
  orx  g0535(.a(n606), .b(n605), .O(n607));
  orx  g0536(.a(n607), .b(n604), .O(n608));
  andx g0537(.a(n590), .b(pi36), .O(n609));
  orx  g0538(.a(n609), .b(pi37), .O(n610));
  andx g0539(.a(n593), .b(pi33), .O(n611));
  andx g0540(.a(n598), .b(pi28), .O(n612));
  orx  g0541(.a(n612), .b(n611), .O(n613));
  andx g0542(.a(n582), .b(pi09), .O(n614));
  andx g0543(.a(n596), .b(pi38), .O(n615));
  orx  g0544(.a(n615), .b(n614), .O(n616));
  orx  g0545(.a(n616), .b(n613), .O(n617));
  orx  g0546(.a(n617), .b(n610), .O(n618));
  orx  g0547(.a(n618), .b(n608), .O(n619));
  andx g0548(.a(n619), .b(n603), .O(n620));
  orx  g0549(.a(n620), .b(n569), .O(n621));
  invx g0550(.a(n558), .O(n622));
  invx g0551(.a(n563), .O(n623));
  andx g0552(.a(n623), .b(n622), .O(n624));
  invx g0553(.a(n624), .O(n625));
  invx g0554(.a(n565), .O(n626));
  andx g0555(.a(n569), .b(n626), .O(n627));
  andx g0556(.a(n627), .b(n304), .O(n628));
  orx  g0557(.a(n628), .b(n625), .O(n629));
  invx g0558(.a(n629), .O(n630));
  andx g0559(.a(n630), .b(n621), .O(n631));
  andx g0560(.a(n631), .b(n567), .O(n632));
  orx  g0561(.a(n632), .b(n564), .O(n633));
  orx  g0562(.a(n633), .b(n561), .O(po00));
  invx g0563(.a(n477), .O(n635));
  andx g0564(.a(n635), .b(pi22), .O(n636));
  andx g0565(.a(n477), .b(n88), .O(n637));
  orx  g0566(.a(n637), .b(n636), .O(n638));
  invx g0567(.a(n638), .O(n639));
  andx g0568(.a(n639), .b(pi33), .O(n640));
  andx g0569(.a(n638), .b(n521), .O(n641));
  orx  g0570(.a(n641), .b(n640), .O(n642));
  invx g0571(.a(n266), .O(n643));
  andx g0572(.a(n643), .b(pi15), .O(n644));
  andx g0573(.a(n266), .b(n223), .O(n645));
  orx  g0574(.a(n645), .b(n644), .O(n646));
  invx g0575(.a(n646), .O(n647));
  andx g0576(.a(n647), .b(pi19), .O(n648));
  andx g0577(.a(n646), .b(n152), .O(n649));
  orx  g0578(.a(n649), .b(n648), .O(n650));
  andx g0579(.a(n650), .b(n642), .O(n651));
  invx g0580(.a(n642), .O(n652));
  invx g0581(.a(n650), .O(n653));
  andx g0582(.a(n653), .b(n652), .O(n654));
  orx  g0583(.a(n654), .b(n651), .O(po01));
  andx g0584(.a(n522), .b(n88), .O(po02));
  orx  g0585(.a(n446), .b(n338), .O(n657));
  andx g0586(.a(n549), .b(n382), .O(n658));
  invx g0587(.a(n658), .O(n659));
  andx g0588(.a(n659), .b(n657), .O(n660));
  invx g0589(.a(n76), .O(n661));
  andx g0590(.a(n547), .b(n661), .O(n662));
  invx g0591(.a(n506), .O(n663));
  andx g0592(.a(n487), .b(n76), .O(n664));
  orx  g0593(.a(n664), .b(n663), .O(n665));
  andx g0594(.a(n665), .b(n501), .O(n666));
  orx  g0595(.a(n666), .b(n662), .O(n667));
  orx  g0596(.a(n667), .b(n660), .O(n668));
  andx g0597(.a(n429), .b(n465), .O(n669));
  orx  g0598(.a(n658), .b(n669), .O(n670));
  invx g0599(.a(n667), .O(n671));
  orx  g0600(.a(n671), .b(n670), .O(n672));
  andx g0601(.a(n672), .b(n668), .O(n673));
  andx g0602(.a(n673), .b(n447), .O(n674));
  andx g0603(.a(n671), .b(n670), .O(n675));
  andx g0604(.a(n667), .b(n660), .O(n676));
  orx  g0605(.a(n676), .b(n675), .O(n677));
  andx g0606(.a(n677), .b(n468), .O(n678));
  orx  g0607(.a(n678), .b(n674), .O(n679));
  andx g0608(.a(n679), .b(n556), .O(n680));
  orx  g0609(.a(n680), .b(n554), .O(n681));
  invx g0610(.a(n662), .O(n682));
  andx g0611(.a(n668), .b(n682), .O(n683));
  andx g0612(.a(n534), .b(n76), .O(n684));
  invx g0613(.a(n684), .O(n685));
  andx g0614(.a(n685), .b(n542), .O(n686));
  andx g0615(.a(n546), .b(n76), .O(n687));
  orx  g0616(.a(n687), .b(n686), .O(n688));
  andx g0617(.a(n671), .b(n468), .O(n689));
  orx  g0618(.a(n689), .b(n688), .O(n690));
  andx g0619(.a(n689), .b(n688), .O(n691));
  invx g0620(.a(n691), .O(n692));
  andx g0621(.a(n692), .b(n690), .O(n693));
  andx g0622(.a(n693), .b(n683), .O(n694));
  orx  g0623(.a(n675), .b(n662), .O(n695));
  invx g0624(.a(n690), .O(n696));
  orx  g0625(.a(n691), .b(n696), .O(n697));
  andx g0626(.a(n697), .b(n695), .O(n698));
  orx  g0627(.a(n698), .b(n694), .O(n699));
  andx g0628(.a(n699), .b(n558), .O(n700));
  andx g0629(.a(n700), .b(n681), .O(n701));
  andx g0630(.a(n699), .b(n563), .O(n702));
  invx g0631(.a(n688), .O(n703));
  andx g0632(.a(n703), .b(n565), .O(n704));
  invx g0633(.a(n569), .O(n705));
  andx g0634(.a(n593), .b(pi26), .O(n706));
  andx g0635(.a(n575), .b(pi16), .O(n707));
  andx g0636(.a(n586), .b(pi18), .O(n708));
  orx  g0637(.a(n708), .b(n707), .O(n709));
  orx  g0638(.a(n709), .b(n706), .O(n710));
  invx g0639(.a(n710), .O(n711));
  andx g0640(.a(n590), .b(pi22), .O(n712));
  invx g0641(.a(n712), .O(n713));
  andx g0642(.a(pi37), .b(n172), .O(n714));
  andx g0643(.a(n714), .b(n713), .O(n715));
  andx g0644(.a(n582), .b(pi13), .O(n716));
  orx  g0645(.a(n716), .b(n612), .O(n717));
  andx g0646(.a(n572), .b(pi15), .O(n718));
  andx g0647(.a(n596), .b(pi19), .O(n719));
  orx  g0648(.a(n719), .b(n718), .O(n720));
  orx  g0649(.a(n720), .b(n717), .O(n721));
  invx g0650(.a(n721), .O(n722));
  andx g0651(.a(n722), .b(n715), .O(n723));
  andx g0652(.a(n723), .b(n711), .O(n724));
  andx g0653(.a(n521), .b(pi27), .O(n725));
  andx g0654(.a(n575), .b(pi09), .O(n726));
  andx g0655(.a(n586), .b(pi47), .O(n727));
  andx g0656(.a(n596), .b(pi41), .O(n728));
  orx  g0657(.a(n728), .b(n727), .O(n729));
  orx  g0658(.a(n729), .b(n726), .O(n730));
  invx g0659(.a(n730), .O(n731));
  andx g0660(.a(n590), .b(pi01), .O(n732));
  invx g0661(.a(n732), .O(n733));
  andx g0662(.a(n95), .b(n172), .O(n734));
  andx g0663(.a(n734), .b(n733), .O(n735));
  andx g0664(.a(n593), .b(pi38), .O(n736));
  andx g0665(.a(n598), .b(pi36), .O(n737));
  orx  g0666(.a(n737), .b(n736), .O(n738));
  andx g0667(.a(n582), .b(pi07), .O(n739));
  andx g0668(.a(n572), .b(pi08), .O(n740));
  orx  g0669(.a(n740), .b(n739), .O(n741));
  orx  g0670(.a(n741), .b(n738), .O(n742));
  invx g0671(.a(n742), .O(n743));
  andx g0672(.a(n743), .b(n735), .O(n744));
  andx g0673(.a(n744), .b(n731), .O(n745));
  orx  g0674(.a(n745), .b(n725), .O(n746));
  orx  g0675(.a(n746), .b(n724), .O(n747));
  andx g0676(.a(n747), .b(n705), .O(n748));
  andx g0677(.a(n627), .b(n521), .O(n749));
  orx  g0678(.a(n749), .b(n625), .O(n750));
  orx  g0679(.a(n750), .b(n748), .O(n751));
  orx  g0680(.a(n751), .b(n704), .O(n752));
  invx g0681(.a(n752), .O(n753));
  orx  g0682(.a(n753), .b(n702), .O(n754));
  orx  g0683(.a(n754), .b(n701), .O(po03));
  andx g0684(.a(n457), .b(n382), .O(n756));
  invx g0685(.a(pi14), .O(n757));
  orx  g0686(.a(n220), .b(n241), .O(n758));
  orx  g0687(.a(n210), .b(n239), .O(n759));
  andx g0688(.a(n759), .b(n758), .O(n760));
  andx g0689(.a(n760), .b(n237), .O(n761));
  orx  g0690(.a(n761), .b(n457), .O(n762));
  andx g0691(.a(n348), .b(n77), .O(n763));
  orx  g0692(.a(n763), .b(n762), .O(n764));
  andx g0693(.a(n457), .b(n77), .O(n765));
  invx g0694(.a(n765), .O(n766));
  andx g0695(.a(n766), .b(n764), .O(n767));
  orx  g0696(.a(n767), .b(n757), .O(n768));
  andx g0697(.a(n362), .b(n77), .O(n769));
  invx g0698(.a(n769), .O(n770));
  andx g0699(.a(n770), .b(n367), .O(n771));
  andx g0700(.a(n769), .b(n453), .O(n772));
  orx  g0701(.a(n772), .b(n771), .O(n773));
  invx g0702(.a(n773), .O(n774));
  orx  g0703(.a(n774), .b(n768), .O(n775));
  invx g0704(.a(n763), .O(n776));
  andx g0705(.a(n776), .b(n353), .O(n777));
  orx  g0706(.a(n765), .b(n777), .O(n778));
  andx g0707(.a(n778), .b(pi14), .O(n779));
  orx  g0708(.a(n773), .b(n779), .O(n780));
  andx g0709(.a(n780), .b(n775), .O(n781));
  andx g0710(.a(n781), .b(n756), .O(n782));
  invx g0711(.a(n756), .O(n783));
  andx g0712(.a(n773), .b(n779), .O(n784));
  andx g0713(.a(n774), .b(n768), .O(n785));
  orx  g0714(.a(n785), .b(n784), .O(n786));
  andx g0715(.a(n786), .b(n783), .O(n787));
  orx  g0716(.a(n787), .b(n782), .O(n788));
  andx g0717(.a(n788), .b(n472), .O(n789));
  invx g0718(.a(n789), .O(n790));
  orx  g0719(.a(n788), .b(n472), .O(n791));
  andx g0720(.a(n791), .b(n558), .O(n792));
  andx g0721(.a(n792), .b(n790), .O(n793));
  orx  g0722(.a(n786), .b(n783), .O(n794));
  orx  g0723(.a(n781), .b(n756), .O(n795));
  andx g0724(.a(n795), .b(n794), .O(n796));
  andx g0725(.a(n796), .b(n563), .O(n797));
  andx g0726(.a(n565), .b(n72), .O(n798));
  andx g0727(.a(n798), .b(n774), .O(n799));
  invx g0728(.a(n799), .O(n800));
  andx g0729(.a(n575), .b(pi33), .O(n801));
  andx g0730(.a(n582), .b(pi38), .O(n802));
  orx  g0731(.a(n802), .b(n712), .O(n803));
  orx  g0732(.a(n803), .b(n801), .O(n804));
  andx g0733(.a(n572), .b(pi36), .O(n805));
  orx  g0734(.a(n805), .b(pi37), .O(n806));
  andx g0735(.a(n598), .b(pi18), .O(n807));
  andx g0736(.a(n586), .b(pi28), .O(n808));
  orx  g0737(.a(n808), .b(n807), .O(n809));
  andx g0738(.a(n596), .b(pi26), .O(n810));
  orx  g0739(.a(n810), .b(n594), .O(n811));
  orx  g0740(.a(n811), .b(n809), .O(n812));
  orx  g0741(.a(n812), .b(n806), .O(n813));
  orx  g0742(.a(n813), .b(n804), .O(n814));
  andx g0743(.a(n586), .b(pi05), .O(n815));
  andx g0744(.a(n572), .b(pi04), .O(n816));
  andx g0745(.a(n593), .b(pi13), .O(n817));
  orx  g0746(.a(n817), .b(n816), .O(n818));
  orx  g0747(.a(n818), .b(n815), .O(n819));
  andx g0748(.a(n590), .b(pi10), .O(n820));
  orx  g0749(.a(n820), .b(n95), .O(n821));
  andx g0750(.a(n596), .b(pi06), .O(n822));
  andx g0751(.a(n598), .b(pi15), .O(n823));
  orx  g0752(.a(n823), .b(n822), .O(n824));
  andx g0753(.a(n575), .b(pi00), .O(n825));
  andx g0754(.a(n582), .b(pi03), .O(n826));
  orx  g0755(.a(n826), .b(n825), .O(n827));
  orx  g0756(.a(n827), .b(n824), .O(n828));
  orx  g0757(.a(n828), .b(n821), .O(n829));
  orx  g0758(.a(n829), .b(n819), .O(n830));
  andx g0759(.a(n830), .b(n814), .O(n831));
  orx  g0760(.a(n831), .b(n569), .O(n832));
  invx g0761(.a(n798), .O(n833));
  andx g0762(.a(n833), .b(n569), .O(n834));
  invx g0763(.a(n834), .O(n835));
  invx g0764(.a(pi21), .O(n836));
  invx g0765(.a(pi25), .O(n837));
  andx g0766(.a(n837), .b(n836), .O(n838));
  andx g0767(.a(pi25), .b(pi21), .O(n839));
  orx  g0768(.a(n839), .b(n838), .O(n840));
  invx g0769(.a(n840), .O(n841));
  invx g0770(.a(pi34), .O(n842));
  andx g0771(.a(n842), .b(pi29), .O(n843));
  andx g0772(.a(pi34), .b(n113), .O(n844));
  orx  g0773(.a(n844), .b(n843), .O(n845));
  invx g0774(.a(n845), .O(n846));
  andx g0775(.a(n846), .b(n841), .O(n847));
  andx g0776(.a(n845), .b(n840), .O(n848));
  orx  g0777(.a(n848), .b(n847), .O(n849));
  invx g0778(.a(n849), .O(n850));
  andx g0779(.a(n850), .b(pi24), .O(n851));
  andx g0780(.a(n302), .b(n223), .O(n852));
  andx g0781(.a(pi26), .b(pi22), .O(n853));
  invx g0782(.a(n853), .O(n854));
  andx g0783(.a(pi28), .b(n176), .O(n855));
  andx g0784(.a(n855), .b(n521), .O(n856));
  andx g0785(.a(n856), .b(n854), .O(n857));
  andx g0786(.a(n857), .b(n852), .O(n858));
  orx  g0787(.a(n858), .b(n148), .O(n859));
  orx  g0788(.a(n859), .b(n851), .O(n860));
  andx g0789(.a(n81), .b(n95), .O(n861));
  invx g0790(.a(n861), .O(n862));
  orx  g0791(.a(n862), .b(n852), .O(n863));
  andx g0792(.a(n147), .b(n136), .O(n864));
  invx g0793(.a(n864), .O(n865));
  andx g0794(.a(n865), .b(n863), .O(n866));
  andx g0795(.a(n866), .b(n860), .O(n867));
  orx  g0796(.a(n867), .b(n835), .O(n868));
  andx g0797(.a(n868), .b(n624), .O(n869));
  andx g0798(.a(n869), .b(n832), .O(n870));
  andx g0799(.a(n870), .b(n800), .O(n871));
  orx  g0800(.a(n871), .b(n797), .O(n872));
  orx  g0801(.a(n872), .b(n793), .O(po04));
  andx g0802(.a(n472), .b(n74), .O(n874));
  orx  g0803(.a(n475), .b(n521), .O(n875));
  invx g0804(.a(n875), .O(n876));
  andx g0805(.a(n876), .b(n558), .O(n877));
  andx g0806(.a(n622), .b(pi43), .O(n878));
  andx g0807(.a(n878), .b(n852), .O(n879));
  orx  g0808(.a(n879), .b(n877), .O(n880));
  orx  g0809(.a(n880), .b(n874), .O(po05));
  andx g0810(.a(n544), .b(n463), .O(n882));
  orx  g0811(.a(n882), .b(n553), .O(po06));
  andx g0812(.a(n337), .b(n326), .O(n884));
  orx  g0813(.a(n884), .b(n465), .O(n885));
  andx g0814(.a(n885), .b(n444), .O(n886));
  invx g0815(.a(n886), .O(n887));
  andx g0816(.a(n445), .b(n625), .O(n888));
  andx g0817(.a(n888), .b(n887), .O(n889));
  andx g0818(.a(n565), .b(n337), .O(n890));
  invx g0819(.a(n890), .O(n891));
  andx g0820(.a(n572), .b(pi06), .O(n892));
  andx g0821(.a(n575), .b(pi10), .O(n893));
  andx g0822(.a(n582), .b(pi05), .O(n894));
  orx  g0823(.a(n894), .b(n893), .O(n895));
  orx  g0824(.a(n895), .b(n892), .O(n896));
  andx g0825(.a(n586), .b(pi13), .O(n897));
  orx  g0826(.a(n897), .b(n95), .O(n898));
  andx g0827(.a(n590), .b(pi16), .O(n899));
  andx g0828(.a(n593), .b(pi18), .O(n900));
  orx  g0829(.a(n900), .b(n899), .O(n901));
  andx g0830(.a(n596), .b(pi15), .O(n902));
  andx g0831(.a(n598), .b(pi19), .O(n903));
  orx  g0832(.a(n903), .b(n902), .O(n904));
  orx  g0833(.a(n904), .b(n901), .O(n905));
  orx  g0834(.a(n905), .b(n898), .O(n906));
  orx  g0835(.a(n906), .b(n896), .O(n907));
  andx g0836(.a(n586), .b(pi38), .O(n908));
  andx g0837(.a(n572), .b(pi41), .O(n909));
  andx g0838(.a(n575), .b(pi01), .O(n910));
  orx  g0839(.a(n910), .b(n909), .O(n911));
  orx  g0840(.a(n911), .b(n908), .O(n912));
  andx g0841(.a(n590), .b(pi33), .O(n913));
  orx  g0842(.a(n913), .b(pi37), .O(n914));
  andx g0843(.a(n593), .b(pi28), .O(n915));
  andx g0844(.a(n598), .b(pi26), .O(n916));
  orx  g0845(.a(n916), .b(n915), .O(n917));
  andx g0846(.a(n582), .b(pi47), .O(n918));
  andx g0847(.a(n596), .b(pi36), .O(n919));
  orx  g0848(.a(n919), .b(n918), .O(n920));
  orx  g0849(.a(n920), .b(n917), .O(n921));
  orx  g0850(.a(n921), .b(n914), .O(n922));
  orx  g0851(.a(n922), .b(n912), .O(n923));
  andx g0852(.a(n923), .b(n907), .O(n924));
  orx  g0853(.a(n924), .b(n569), .O(n925));
  andx g0854(.a(n627), .b(n88), .O(n926));
  orx  g0855(.a(n926), .b(n625), .O(n927));
  invx g0856(.a(n927), .O(n928));
  andx g0857(.a(n928), .b(n925), .O(n929));
  andx g0858(.a(n929), .b(n891), .O(n930));
  orx  g0859(.a(n930), .b(n889), .O(po07));
  andx g0860(.a(n370), .b(n77), .O(n932));
  orx  g0861(.a(n932), .b(n435), .O(n933));
  andx g0862(.a(n434), .b(n77), .O(n934));
  invx g0863(.a(n934), .O(n935));
  andx g0864(.a(n935), .b(n933), .O(n936));
  andx g0865(.a(n936), .b(n798), .O(n937));
  invx g0866(.a(n937), .O(n938));
  andx g0867(.a(n575), .b(pi38), .O(n939));
  andx g0868(.a(n596), .b(pi33), .O(n940));
  orx  g0869(.a(n940), .b(n599), .O(n941));
  orx  g0870(.a(n941), .b(n939), .O(n942));
  andx g0871(.a(n572), .b(pi01), .O(n943));
  orx  g0872(.a(n943), .b(pi37), .O(n944));
  andx g0873(.a(n582), .b(pi41), .O(n945));
  andx g0874(.a(n586), .b(pi36), .O(n946));
  orx  g0875(.a(n946), .b(n945), .O(n947));
  andx g0876(.a(n590), .b(pi28), .O(n948));
  orx  g0877(.a(n948), .b(n706), .O(n949));
  orx  g0878(.a(n949), .b(n947), .O(n950));
  orx  g0879(.a(n950), .b(n944), .O(n951));
  orx  g0880(.a(n951), .b(n942), .O(n952));
  andx g0881(.a(n590), .b(pi15), .O(n953));
  andx g0882(.a(n582), .b(pi00), .O(n954));
  andx g0883(.a(n575), .b(pi06), .O(n955));
  orx  g0884(.a(n955), .b(n954), .O(n956));
  orx  g0885(.a(n956), .b(n953), .O(n957));
  andx g0886(.a(n572), .b(pi05), .O(n958));
  orx  g0887(.a(n958), .b(n95), .O(n959));
  andx g0888(.a(n593), .b(pi16), .O(n960));
  andx g0889(.a(n586), .b(pi10), .O(n961));
  orx  g0890(.a(n961), .b(n960), .O(n962));
  andx g0891(.a(n596), .b(pi13), .O(n963));
  orx  g0892(.a(n963), .b(n807), .O(n964));
  orx  g0893(.a(n964), .b(n962), .O(n965));
  orx  g0894(.a(n965), .b(n959), .O(n966));
  orx  g0895(.a(n966), .b(n957), .O(n967));
  andx g0896(.a(n967), .b(n952), .O(n968));
  orx  g0897(.a(n968), .b(n569), .O(n969));
  andx g0898(.a(n217), .b(n180), .O(n970));
  andx g0899(.a(pi12), .b(pi11), .O(n971));
  orx  g0900(.a(n971), .b(n970), .O(n972));
  invx g0901(.a(n972), .O(n973));
  andx g0902(.a(n162), .b(pi20), .O(n974));
  andx g0903(.a(pi17), .b(n160), .O(n975));
  orx  g0904(.a(n975), .b(n974), .O(n976));
  invx g0905(.a(n976), .O(n977));
  andx g0906(.a(n977), .b(n973), .O(n978));
  andx g0907(.a(n976), .b(n972), .O(n979));
  orx  g0908(.a(n979), .b(n978), .O(n980));
  invx g0909(.a(n980), .O(n981));
  andx g0910(.a(n981), .b(n82), .O(n982));
  andx g0911(.a(n147), .b(pi19), .O(n983));
  orx  g0912(.a(n983), .b(n835), .O(n984));
  orx  g0913(.a(n984), .b(n982), .O(n985));
  andx g0914(.a(n985), .b(n624), .O(n986));
  andx g0915(.a(n986), .b(n969), .O(n987));
  andx g0916(.a(n987), .b(n938), .O(n988));
  andx g0917(.a(n444), .b(n326), .O(n989));
  andx g0918(.a(n796), .b(n989), .O(n990));
  andx g0919(.a(n773), .b(n457), .O(n991));
  orx  g0920(.a(n991), .b(n454), .O(n992));
  andx g0921(.a(n992), .b(n382), .O(n993));
  invx g0922(.a(n993), .O(n994));
  andx g0923(.a(n271), .b(n77), .O(n995));
  orx  g0924(.a(n995), .b(n439), .O(n996));
  andx g0925(.a(n438), .b(n77), .O(n997));
  invx g0926(.a(n997), .O(n998));
  andx g0927(.a(n998), .b(n996), .O(n999));
  invx g0928(.a(n999), .O(n1000));
  andx g0929(.a(n1000), .b(n784), .O(n1001));
  andx g0930(.a(n999), .b(n775), .O(n1002));
  orx  g0931(.a(n1002), .b(n1001), .O(n1003));
  orx  g0932(.a(n1003), .b(n994), .O(n1004));
  orx  g0933(.a(n999), .b(n775), .O(n1005));
  orx  g0934(.a(n1000), .b(n784), .O(n1006));
  andx g0935(.a(n1006), .b(n1005), .O(n1007));
  orx  g0936(.a(n1007), .b(n993), .O(n1008));
  andx g0937(.a(n1008), .b(n1004), .O(n1009));
  andx g0938(.a(n1009), .b(n990), .O(n1010));
  orx  g0939(.a(n1010), .b(n472), .O(n1011));
  andx g0940(.a(n1011), .b(n558), .O(n1012));
  orx  g0941(.a(n1012), .b(n563), .O(n1013));
  andx g0942(.a(n461), .b(n382), .O(n1014));
  invx g0943(.a(n1014), .O(n1015));
  andx g0944(.a(n1005), .b(n1015), .O(n1016));
  andx g0945(.a(n1016), .b(n936), .O(n1017));
  invx g0946(.a(n1017), .O(n1018));
  orx  g0947(.a(n1016), .b(n936), .O(n1019));
  andx g0948(.a(n1019), .b(n1018), .O(n1020));
  andx g0949(.a(n1020), .b(n1013), .O(n1021));
  orx  g0950(.a(n1021), .b(n988), .O(po08));
  andx g0951(.a(n981), .b(n850), .O(n1023));
  andx g0952(.a(n980), .b(n849), .O(n1024));
  orx  g0953(.a(n1024), .b(n1023), .O(po09));
  invx g0954(.a(n264), .O(n1026));
  andx g0955(.a(n1026), .b(pi19), .O(n1027));
  invx g0956(.a(n1027), .O(po10));
  orx  g0957(.a(n993), .b(n784), .O(po11));
  orx  g0958(.a(n677), .b(n468), .O(n1030));
  orx  g0959(.a(n673), .b(n447), .O(n1031));
  andx g0960(.a(n1031), .b(n1030), .O(n1032));
  orx  g0961(.a(n1032), .b(n557), .O(n1033));
  andx g0962(.a(n1033), .b(n555), .O(n1034));
  orx  g0963(.a(n697), .b(n695), .O(n1035));
  orx  g0964(.a(n693), .b(n683), .O(n1036));
  andx g0965(.a(n1036), .b(n1035), .O(n1037));
  orx  g0966(.a(n1037), .b(n622), .O(n1038));
  orx  g0967(.a(n1038), .b(n1034), .O(n1039));
  orx  g0968(.a(n1037), .b(n623), .O(n1040));
  andx g0969(.a(n752), .b(n1040), .O(n1041));
  andx g0970(.a(n1041), .b(n1039), .O(n1042));
  andx g0971(.a(n1032), .b(n557), .O(n1043));
  orx  g0972(.a(n1043), .b(n622), .O(n1044));
  orx  g0973(.a(n1044), .b(n680), .O(n1045));
  orx  g0974(.a(n1032), .b(n623), .O(n1046));
  andx g0975(.a(n667), .b(n565), .O(n1047));
  invx g0976(.a(n1047), .O(n1048));
  andx g0977(.a(n582), .b(pi10), .O(n1049));
  andx g0978(.a(n575), .b(pi15), .O(n1050));
  orx  g0979(.a(n1050), .b(n916), .O(n1051));
  orx  g0980(.a(n1051), .b(n1049), .O(n1052));
  andx g0981(.a(n586), .b(pi16), .O(n1053));
  orx  g0982(.a(n1053), .b(n95), .O(n1054));
  andx g0983(.a(n572), .b(pi13), .O(n1055));
  andx g0984(.a(n593), .b(pi22), .O(n1056));
  orx  g0985(.a(n1056), .b(n1055), .O(n1057));
  andx g0986(.a(n596), .b(pi18), .O(n1058));
  andx g0987(.a(n590), .b(pi19), .O(n1059));
  orx  g0988(.a(n1059), .b(n1058), .O(n1060));
  orx  g0989(.a(n1060), .b(n1057), .O(n1061));
  orx  g0990(.a(n1061), .b(n1054), .O(n1062));
  orx  g0991(.a(n1062), .b(n1052), .O(n1063));
  andx g0992(.a(n586), .b(pi41), .O(n1064));
  andx g0993(.a(n572), .b(pi09), .O(n1065));
  andx g0994(.a(n575), .b(pi47), .O(n1066));
  orx  g0995(.a(n1066), .b(n1065), .O(n1067));
  orx  g0996(.a(n1067), .b(n1064), .O(n1068));
  andx g0997(.a(n590), .b(pi38), .O(n1069));
  orx  g0998(.a(n1069), .b(pi37), .O(n1070));
  andx g0999(.a(n593), .b(pi36), .O(n1071));
  andx g1000(.a(n598), .b(pi33), .O(n1072));
  orx  g1001(.a(n1072), .b(n1071), .O(n1073));
  andx g1002(.a(n582), .b(pi08), .O(n1074));
  andx g1003(.a(n596), .b(pi01), .O(n1075));
  orx  g1004(.a(n1075), .b(n1074), .O(n1076));
  orx  g1005(.a(n1076), .b(n1073), .O(n1077));
  orx  g1006(.a(n1077), .b(n1070), .O(n1078));
  orx  g1007(.a(n1078), .b(n1068), .O(n1079));
  andx g1008(.a(n1079), .b(n1063), .O(n1080));
  orx  g1009(.a(n1080), .b(n569), .O(n1081));
  andx g1010(.a(n627), .b(n474), .O(n1082));
  orx  g1011(.a(n1082), .b(n625), .O(n1083));
  invx g1012(.a(n1083), .O(n1084));
  andx g1013(.a(n1084), .b(n1081), .O(n1085));
  andx g1014(.a(n1085), .b(n1048), .O(n1086));
  invx g1015(.a(n1086), .O(n1087));
  andx g1016(.a(n1087), .b(n1046), .O(n1088));
  andx g1017(.a(n1088), .b(n1045), .O(n1089));
  orx  g1018(.a(n1089), .b(n1042), .O(n1090));
  orx  g1019(.a(n679), .b(n556), .O(n1091));
  andx g1020(.a(n1091), .b(n558), .O(n1092));
  andx g1021(.a(n1092), .b(n1033), .O(n1093));
  andx g1022(.a(n679), .b(n563), .O(n1094));
  orx  g1023(.a(n1086), .b(n1094), .O(n1095));
  orx  g1024(.a(n1095), .b(n1093), .O(po17));
  orx  g1025(.a(po17), .b(po03), .O(n1097));
  andx g1026(.a(n1097), .b(n1090), .O(n1098));
  andx g1027(.a(n1007), .b(n993), .O(n1099));
  andx g1028(.a(n1003), .b(n994), .O(n1100));
  orx  g1029(.a(n1100), .b(n1099), .O(n1101));
  andx g1030(.a(n1101), .b(n791), .O(n1102));
  orx  g1031(.a(n1102), .b(n622), .O(n1103));
  orx  g1032(.a(n1103), .b(n1010), .O(n1104));
  andx g1033(.a(n1009), .b(n563), .O(n1105));
  andx g1034(.a(n999), .b(n798), .O(n1106));
  invx g1035(.a(n1106), .O(n1107));
  andx g1036(.a(n575), .b(pi36), .O(n1108));
  andx g1037(.a(n596), .b(pi28), .O(n1109));
  orx  g1038(.a(n1109), .b(n1056), .O(n1110));
  orx  g1039(.a(n1110), .b(n1108), .O(n1111));
  andx g1040(.a(n572), .b(pi38), .O(n1112));
  orx  g1041(.a(n1112), .b(pi37), .O(n1113));
  andx g1042(.a(n582), .b(pi01), .O(n1114));
  andx g1043(.a(n586), .b(pi33), .O(n1115));
  orx  g1044(.a(n1115), .b(n1114), .O(n1116));
  andx g1045(.a(n590), .b(pi26), .O(n1117));
  orx  g1046(.a(n1117), .b(n903), .O(n1118));
  orx  g1047(.a(n1118), .b(n1116), .O(n1119));
  orx  g1048(.a(n1119), .b(n1113), .O(n1120));
  orx  g1049(.a(n1120), .b(n1111), .O(n1121));
  andx g1050(.a(n586), .b(pi06), .O(n1122));
  andx g1051(.a(n572), .b(pi00), .O(n1123));
  andx g1052(.a(n593), .b(pi15), .O(n1124));
  orx  g1053(.a(n1124), .b(n1123), .O(n1125));
  orx  g1054(.a(n1125), .b(n1122), .O(n1126));
  andx g1055(.a(n590), .b(pi13), .O(n1127));
  orx  g1056(.a(n1127), .b(n95), .O(n1128));
  andx g1057(.a(n596), .b(pi10), .O(n1129));
  andx g1058(.a(n598), .b(pi16), .O(n1130));
  orx  g1059(.a(n1130), .b(n1129), .O(n1131));
  andx g1060(.a(n575), .b(pi05), .O(n1132));
  andx g1061(.a(n582), .b(pi04), .O(n1133));
  orx  g1062(.a(n1133), .b(n1132), .O(n1134));
  orx  g1063(.a(n1134), .b(n1131), .O(n1135));
  orx  g1064(.a(n1135), .b(n1128), .O(n1136));
  orx  g1065(.a(n1136), .b(n1126), .O(n1137));
  andx g1066(.a(n1137), .b(n1121), .O(n1138));
  orx  g1067(.a(n1138), .b(n569), .O(n1139));
  andx g1068(.a(n650), .b(n82), .O(n1140));
  andx g1069(.a(n147), .b(pi18), .O(n1141));
  orx  g1070(.a(n1141), .b(n835), .O(n1142));
  orx  g1071(.a(n1142), .b(n1140), .O(n1143));
  andx g1072(.a(n1143), .b(n624), .O(n1144));
  andx g1073(.a(n1144), .b(n1139), .O(n1145));
  andx g1074(.a(n1145), .b(n1107), .O(n1146));
  orx  g1075(.a(n1146), .b(n1105), .O(n1147));
  invx g1076(.a(n1147), .O(n1148));
  andx g1077(.a(n1148), .b(n1104), .O(n1149));
  invx g1078(.a(n1149), .O(po18));
  andx g1079(.a(po18), .b(po08), .O(n1151));
  invx g1080(.a(n988), .O(n1152));
  orx  g1081(.a(n1101), .b(n791), .O(n1153));
  andx g1082(.a(n1153), .b(n989), .O(n1154));
  orx  g1083(.a(n1154), .b(n622), .O(n1155));
  andx g1084(.a(n1155), .b(n623), .O(n1156));
  invx g1085(.a(n1020), .O(n1157));
  orx  g1086(.a(n1157), .b(n1156), .O(n1158));
  andx g1087(.a(n1158), .b(n1152), .O(n1159));
  andx g1088(.a(n1149), .b(n1159), .O(n1160));
  orx  g1089(.a(n1160), .b(n1151), .O(n1161));
  andx g1090(.a(n798), .b(n767), .O(n1162));
  invx g1091(.a(n1162), .O(n1163));
  andx g1092(.a(n642), .b(pi24), .O(n1164));
  andx g1093(.a(n876), .b(n176), .O(n1165));
  orx  g1094(.a(n1165), .b(n148), .O(n1166));
  orx  g1095(.a(n1166), .b(n1164), .O(n1167));
  andx g1096(.a(po10), .b(n861), .O(n1168));
  andx g1097(.a(n147), .b(n223), .O(n1169));
  orx  g1098(.a(n1169), .b(n1168), .O(n1170));
  invx g1099(.a(n1170), .O(n1171));
  andx g1100(.a(n1171), .b(n1167), .O(n1172));
  orx  g1101(.a(n1172), .b(n835), .O(n1173));
  andx g1102(.a(n575), .b(pi28), .O(n1174));
  andx g1103(.a(n596), .b(pi22), .O(n1175));
  orx  g1104(.a(n1175), .b(n1059), .O(n1176));
  orx  g1105(.a(n1176), .b(n1174), .O(n1177));
  andx g1106(.a(n572), .b(pi33), .O(n1178));
  orx  g1107(.a(n1178), .b(pi37), .O(n1179));
  andx g1108(.a(n582), .b(pi36), .O(n1180));
  orx  g1109(.a(n1180), .b(n1130), .O(n1181));
  andx g1110(.a(n586), .b(pi26), .O(n1182));
  orx  g1111(.a(n1182), .b(n900), .O(n1183));
  orx  g1112(.a(n1183), .b(n1181), .O(n1184));
  orx  g1113(.a(n1184), .b(n1179), .O(n1185));
  orx  g1114(.a(n1185), .b(n1177), .O(n1186));
  andx g1115(.a(n586), .b(pi00), .O(n1187));
  andx g1116(.a(n572), .b(pi03), .O(n1188));
  andx g1117(.a(n593), .b(pi10), .O(n1189));
  orx  g1118(.a(n1189), .b(n1188), .O(n1190));
  orx  g1119(.a(n1190), .b(n1187), .O(n1191));
  andx g1120(.a(n590), .b(pi06), .O(n1192));
  orx  g1121(.a(n1192), .b(n95), .O(n1193));
  andx g1122(.a(n596), .b(pi05), .O(n1194));
  andx g1123(.a(n598), .b(pi13), .O(n1195));
  orx  g1124(.a(n1195), .b(n1194), .O(n1196));
  andx g1125(.a(n575), .b(pi04), .O(n1197));
  andx g1126(.a(n582), .b(pi02), .O(n1198));
  orx  g1127(.a(n1198), .b(n1197), .O(n1199));
  orx  g1128(.a(n1199), .b(n1196), .O(n1200));
  orx  g1129(.a(n1200), .b(n1193), .O(n1201));
  orx  g1130(.a(n1201), .b(n1191), .O(n1202));
  andx g1131(.a(n1202), .b(n1186), .O(n1203));
  orx  g1132(.a(n1203), .b(n569), .O(n1204));
  andx g1133(.a(n1204), .b(n624), .O(n1205));
  andx g1134(.a(n1205), .b(n1173), .O(n1206));
  andx g1135(.a(n1206), .b(n1163), .O(n1207));
  andx g1136(.a(n767), .b(n757), .O(n1208));
  invx g1137(.a(n1208), .O(n1209));
  andx g1138(.a(n768), .b(n625), .O(n1210));
  andx g1139(.a(n1210), .b(n1209), .O(n1211));
  orx  g1140(.a(n1211), .b(n1207), .O(po14));
  invx g1141(.a(po14), .O(n1213));
  andx g1142(.a(n1213), .b(n1161), .O(n1214));
  orx  g1143(.a(n1149), .b(n1159), .O(n1215));
  orx  g1144(.a(po18), .b(po08), .O(n1216));
  andx g1145(.a(n1216), .b(n1215), .O(n1217));
  andx g1146(.a(po14), .b(n1217), .O(n1218));
  orx  g1147(.a(n1218), .b(n1214), .O(n1219));
  orx  g1148(.a(n469), .b(n466), .O(n1220));
  orx  g1149(.a(n448), .b(n339), .O(n1221));
  andx g1150(.a(n1221), .b(n1220), .O(n1222));
  andx g1151(.a(n554), .b(n1222), .O(n1223));
  orx  g1152(.a(n1223), .b(n622), .O(n1224));
  orx  g1153(.a(n1224), .b(n556), .O(n1225));
  invx g1154(.a(n633), .O(n1226));
  andx g1155(.a(n1226), .b(n1225), .O(n1227));
  invx g1156(.a(po07), .O(n1228));
  orx  g1157(.a(n1228), .b(n1227), .O(n1229));
  orx  g1158(.a(po07), .b(po00), .O(n1230));
  andx g1159(.a(n1230), .b(n1229), .O(n1231));
  andx g1160(.a(n1231), .b(po04), .O(n1232));
  invx g1161(.a(po04), .O(n1233));
  andx g1162(.a(po07), .b(po00), .O(n1234));
  andx g1163(.a(n1228), .b(n1227), .O(n1235));
  orx  g1164(.a(n1235), .b(n1234), .O(n1236));
  andx g1165(.a(n1236), .b(n1233), .O(n1237));
  orx  g1166(.a(n1237), .b(n1232), .O(n1238));
  orx  g1167(.a(n1238), .b(n1219), .O(n1239));
  orx  g1168(.a(po14), .b(n1217), .O(n1240));
  orx  g1169(.a(n1213), .b(n1161), .O(n1241));
  andx g1170(.a(n1241), .b(n1240), .O(n1242));
  orx  g1171(.a(n1236), .b(n1233), .O(n1243));
  orx  g1172(.a(n1231), .b(po04), .O(n1244));
  andx g1173(.a(n1244), .b(n1243), .O(n1245));
  orx  g1174(.a(n1245), .b(n1242), .O(n1246));
  andx g1175(.a(n1246), .b(n1239), .O(n1247));
  andx g1176(.a(n1247), .b(n1098), .O(n1248));
  andx g1177(.a(po17), .b(po03), .O(n1249));
  andx g1178(.a(n1089), .b(n1042), .O(n1250));
  orx  g1179(.a(n1250), .b(n1249), .O(n1251));
  andx g1180(.a(n1245), .b(n1242), .O(n1252));
  andx g1181(.a(n1238), .b(n1219), .O(n1253));
  orx  g1182(.a(n1253), .b(n1252), .O(n1254));
  andx g1183(.a(n1254), .b(n1251), .O(n1255));
  orx  g1184(.a(n1255), .b(n1248), .O(po12));
  andx g1185(.a(n544), .b(n376), .O(po13));
  invx g1186(.a(pi45), .O(n1258));
  orx  g1187(.a(n1258), .b(pi46), .O(n1259));
  invx g1188(.a(n1259), .O(n1260));
  orx  g1189(.a(n1260), .b(n1098), .O(n1261));
  orx  g1190(.a(n1259), .b(pi49), .O(n1262));
  andx g1191(.a(n1262), .b(n1261), .O(n1263));
  orx  g1192(.a(n1263), .b(n1254), .O(n1264));
  andx g1193(.a(n1259), .b(n1251), .O(n1265));
  invx g1194(.a(n1262), .O(n1266));
  orx  g1195(.a(n1266), .b(n1265), .O(n1267));
  orx  g1196(.a(n1267), .b(n1247), .O(n1268));
  andx g1197(.a(n1268), .b(n1264), .O(po15));
  andx g1198(.a(n1213), .b(n1233), .O(n1270));
  andx g1199(.a(n1270), .b(n1235), .O(n1271));
  andx g1200(.a(n1271), .b(n1160), .O(n1272));
  andx g1201(.a(n1272), .b(n1250), .O(n1273));
  andx g1202(.a(n1260), .b(n1250), .O(n1274));
  orx  g1203(.a(n1274), .b(n1258), .O(n1275));
  orx  g1204(.a(n1275), .b(n1273), .O(po16));
  andx g1205(.a(pi43), .b(pi40), .O(n1277));
  orx  g1206(.a(n152), .b(n160), .O(n1278));
  orx  g1207(.a(n180), .b(n136), .O(n1279));
  andx g1208(.a(n1279), .b(n1278), .O(n1280));
  orx  g1209(.a(n113), .b(n474), .O(n1281));
  orx  g1210(.a(n230), .b(n162), .O(n1282));
  andx g1211(.a(n1282), .b(n1281), .O(n1283));
  andx g1212(.a(n1283), .b(n1280), .O(n1284));
  orx  g1213(.a(n217), .b(n223), .O(n1285));
  orx  g1214(.a(n88), .b(n836), .O(n1286));
  andx g1215(.a(n1286), .b(n1285), .O(n1287));
  orx  g1216(.a(n842), .b(n521), .O(n1288));
  orx  g1217(.a(n304), .b(n837), .O(n1289));
  andx g1218(.a(n1289), .b(n1288), .O(n1290));
  andx g1219(.a(n1290), .b(n1287), .O(n1291));
  andx g1220(.a(n1291), .b(n1284), .O(n1292));
  orx  g1221(.a(n1292), .b(n1277), .O(n1293));
  andx g1222(.a(n89), .b(pi43), .O(n1294));
  invx g1223(.a(n1294), .O(n1295));
  orx  g1224(.a(n1295), .b(n875), .O(n1296));
  andx g1225(.a(n180), .b(n162), .O(n1297));
  orx  g1226(.a(n1297), .b(n160), .O(n1298));
  orx  g1227(.a(n1298), .b(n147), .O(n1299));
  andx g1228(.a(n1299), .b(n1296), .O(n1300));
  andx g1229(.a(n1300), .b(n1293), .O(po19));
  andx g1230(.a(n544), .b(n464), .O(n1302));
  orx  g1231(.a(n1302), .b(n553), .O(n1303));
  invx g1232(.a(n544), .O(n1304));
  andx g1233(.a(n429), .b(n336), .O(n1305));
  andx g1234(.a(n1305), .b(n671), .O(n1306));
  invx g1235(.a(n1306), .O(n1307));
  andx g1236(.a(n1307), .b(n1304), .O(n1308));
  andx g1237(.a(n1306), .b(n544), .O(n1309));
  orx  g1238(.a(n1309), .b(n444), .O(n1310));
  orx  g1239(.a(n1310), .b(n1308), .O(n1311));
  invx g1240(.a(n1311), .O(n1312));
  andx g1241(.a(n1312), .b(n1303), .O(n1313));
  invx g1242(.a(n1313), .O(n1314));
  orx  g1243(.a(n1312), .b(n1303), .O(n1315));
  andx g1244(.a(n1315), .b(n1314), .O(n1316));
  invx g1245(.a(n1316), .O(n1317));
  orx  g1246(.a(n1317), .b(n683), .O(n1318));
  orx  g1247(.a(n1316), .b(n695), .O(n1319));
  andx g1248(.a(n1295), .b(n146), .O(n1320));
  andx g1249(.a(n1320), .b(n1319), .O(n1321));
  andx g1250(.a(n1321), .b(n1318), .O(n1322));
  andx g1251(.a(n1294), .b(n644), .O(n1323));
  orx  g1252(.a(n636), .b(n521), .O(n1324));
  orx  g1253(.a(pi33), .b(pi26), .O(n1325));
  andx g1254(.a(n1325), .b(n80), .O(n1326));
  andx g1255(.a(n1326), .b(n1324), .O(n1327));
  orx  g1256(.a(n1327), .b(n1323), .O(n1328));
  orx  g1257(.a(n1328), .b(n1322), .O(po20));
  invx g1258(.a(n1273), .O(po21));
endmodule


