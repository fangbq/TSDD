// Benchmark "top" written by ABC on Fri Feb  7 13:31:43 2014

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122;
  wire n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n456, n457, n458,
    n459, n460, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1217, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1298,
    n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1496, n1497, n1498, n1499, n1500, n1501,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1521, n1522, n1523, n1524, n1525,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1540, n1541, n1542, n1543, n1544, n1545, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1578, n1579, n1580, n1581,
    n1582, n1583, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1605, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1615, n1618,
    n1619, n1620, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1674,
    n1675, n1676, n1677, n1678, n1679, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
    n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1758,
    n1759, n1760, n1761, n1762, n1763, n1765, n1766, n1767, n1768, n1770,
    n1771, n1772, n1775, n1776, n1777, n1778, n1779, n1780, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1793, n1794, n1795, n1796, n1797,
    n1798, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1816, n1817, n1818, n1819, n1821,
    n1822, n1823, n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832,
    n1833, n1836, n1837, n1838, n1839, n1840, n1841, n1845, n1846, n1847,
    n1848, n1849, n1850, n1853, n1854, n1855, n1856, n1858, n1859, n1860,
    n1861, n1862, n1863, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
    n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1901, n1902,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1912, n1913, n1914,
    n1915, n1916, n1917, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1929, n1930, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1946, n1947, n1948, n1949, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1959, n1961, n1962, n1963, n1964,
    n1965, n1966;
  invx g0000(.a(pi023), .O(n301));
  invx g0001(.a(pi022), .O(n302));
  andx g0002(.a(n302), .b(pi028), .O(n303));
  orx  g0003(.a(pi024), .b(pi028), .O(n304));
  invx g0004(.a(n304), .O(n305));
  orx  g0005(.a(n305), .b(n303), .O(n306));
  orx  g0006(.a(n306), .b(n301), .O(n307));
  invx g0007(.a(pi026), .O(n308));
  invx g0008(.a(pi025), .O(n309));
  andx g0009(.a(n309), .b(pi028), .O(n310));
  invx g0010(.a(pi028), .O(n311));
  invx g0011(.a(pi027), .O(n312));
  andx g0012(.a(n312), .b(n311), .O(n313));
  orx  g0013(.a(n313), .b(n310), .O(n314));
  orx  g0014(.a(n314), .b(n308), .O(n315));
  andx g0015(.a(n315), .b(n307), .O(n316));
  orx  g0016(.a(pi025), .b(n311), .O(n317));
  orx  g0017(.a(pi027), .b(pi028), .O(n318));
  andx g0018(.a(n318), .b(n317), .O(n319));
  andx g0019(.a(n319), .b(pi026), .O(n320));
  andx g0020(.a(n314), .b(n308), .O(n321));
  orx  g0021(.a(n321), .b(n320), .O(n322));
  invx g0022(.a(pi031), .O(n323));
  invx g0023(.a(pi029), .O(n324));
  andx g0024(.a(n324), .b(pi028), .O(n325));
  orx  g0025(.a(pi030), .b(pi028), .O(n326));
  invx g0026(.a(n326), .O(n327));
  orx  g0027(.a(n327), .b(n325), .O(n328));
  orx  g0028(.a(n328), .b(n323), .O(n329));
  orx  g0029(.a(n329), .b(n322), .O(n330));
  andx g0030(.a(n330), .b(n316), .O(n331));
  andx g0031(.a(n306), .b(n301), .O(n332));
  orx  g0032(.a(n332), .b(n331), .O(n333));
  orx  g0033(.a(pi019), .b(n311), .O(n334));
  invx g0034(.a(pi021), .O(n335));
  andx g0035(.a(n335), .b(n311), .O(n336));
  invx g0036(.a(n336), .O(n337));
  andx g0037(.a(n337), .b(n334), .O(n338));
  andx g0038(.a(n338), .b(pi020), .O(n339));
  invx g0039(.a(n339), .O(n340));
  andx g0040(.a(n340), .b(n333), .O(n341));
  orx  g0041(.a(n338), .b(pi020), .O(n342));
  invx g0042(.a(n342), .O(n343));
  orx  g0043(.a(n343), .b(n341), .O(n344));
  orx  g0044(.a(pi016), .b(n311), .O(n345));
  invx g0045(.a(pi018), .O(n346));
  andx g0046(.a(n346), .b(n311), .O(n347));
  invx g0047(.a(n347), .O(n348));
  andx g0048(.a(n348), .b(n345), .O(n349));
  andx g0049(.a(n349), .b(pi017), .O(n350));
  invx g0050(.a(n350), .O(n351));
  andx g0051(.a(n351), .b(n344), .O(n352));
  invx g0052(.a(pi017), .O(n353));
  invx g0053(.a(n349), .O(n354));
  andx g0054(.a(n354), .b(n353), .O(n355));
  orx  g0055(.a(n355), .b(n352), .O(n356));
  invx g0056(.a(n356), .O(n357));
  orx  g0057(.a(pi000), .b(n311), .O(n358));
  invx g0058(.a(pi009), .O(n359));
  andx g0059(.a(n359), .b(n311), .O(n360));
  invx g0060(.a(n360), .O(n361));
  andx g0061(.a(n361), .b(n358), .O(n362));
  andx g0062(.a(n362), .b(pi010), .O(n363));
  invx g0063(.a(pi010), .O(n364));
  invx g0064(.a(n362), .O(n365));
  andx g0065(.a(n365), .b(n364), .O(n366));
  orx  g0066(.a(n366), .b(n363), .O(n367));
  invx g0067(.a(n367), .O(n368));
  orx  g0068(.a(pi008), .b(n311), .O(n369));
  invx g0069(.a(pi012), .O(n370));
  andx g0070(.a(n370), .b(n311), .O(n371));
  invx g0071(.a(n371), .O(n372));
  andx g0072(.a(n372), .b(n369), .O(n373));
  andx g0073(.a(n373), .b(pi011), .O(n374));
  invx g0074(.a(n374), .O(n375));
  invx g0075(.a(pi011), .O(n376));
  invx g0076(.a(n373), .O(n377));
  andx g0077(.a(n377), .b(n376), .O(n378));
  invx g0078(.a(n378), .O(n379));
  andx g0079(.a(n379), .b(n375), .O(n380));
  invx g0080(.a(pi014), .O(n381));
  orx  g0081(.a(pi013), .b(n311), .O(n382));
  invx g0082(.a(pi015), .O(n383));
  andx g0083(.a(n383), .b(n311), .O(n384));
  invx g0084(.a(n384), .O(n385));
  andx g0085(.a(n385), .b(n382), .O(n386));
  invx g0086(.a(n386), .O(n387));
  andx g0087(.a(n387), .b(n381), .O(n388));
  invx g0088(.a(n388), .O(n389));
  andx g0089(.a(n386), .b(pi014), .O(n390));
  invx g0090(.a(n390), .O(n391));
  andx g0091(.a(n391), .b(n389), .O(n392));
  andx g0092(.a(n392), .b(n380), .O(n393));
  andx g0093(.a(n393), .b(n368), .O(n394));
  invx g0094(.a(pi037), .O(n395));
  orx  g0095(.a(pi035), .b(n311), .O(n396));
  invx g0096(.a(pi036), .O(n397));
  andx g0097(.a(n397), .b(n311), .O(n398));
  invx g0098(.a(n398), .O(n399));
  andx g0099(.a(n399), .b(n396), .O(n400));
  invx g0100(.a(n400), .O(n401));
  andx g0101(.a(n401), .b(n395), .O(n402));
  andx g0102(.a(n400), .b(pi037), .O(n403));
  orx  g0103(.a(n403), .b(n402), .O(n404));
  invx g0104(.a(n404), .O(n405));
  andx g0105(.a(n405), .b(n394), .O(n406));
  andx g0106(.a(n406), .b(n357), .O(n407));
  invx g0107(.a(n402), .O(n408));
  invx g0108(.a(n363), .O(n409));
  orx  g0109(.a(n375), .b(n367), .O(n410));
  andx g0110(.a(n410), .b(n409), .O(n411));
  orx  g0111(.a(n411), .b(n388), .O(n412));
  andx g0112(.a(n412), .b(n391), .O(n413));
  invx g0113(.a(n413), .O(n414));
  andx g0114(.a(n414), .b(n408), .O(n415));
  orx  g0115(.a(n415), .b(n403), .O(n416));
  orx  g0116(.a(n416), .b(n407), .O(po000));
  invx g0117(.a(pi177), .O(po001));
  invx g0118(.a(pi079), .O(n419));
  andx g0119(.a(pi064), .b(n419), .O(n420));
  invx g0120(.a(n420), .O(n421));
  orx  g0121(.a(pi029), .b(n311), .O(n422));
  andx g0122(.a(n326), .b(n422), .O(n423));
  andx g0123(.a(n423), .b(pi031), .O(n424));
  andx g0124(.a(n328), .b(n323), .O(n425));
  orx  g0125(.a(n425), .b(n424), .O(n426));
  invx g0126(.a(n426), .O(n427));
  andx g0127(.a(n427), .b(pi032), .O(n428));
  invx g0128(.a(n428), .O(n429));
  andx g0129(.a(n429), .b(n329), .O(n430));
  andx g0130(.a(n430), .b(n322), .O(n431));
  orx  g0131(.a(n430), .b(n322), .O(n432));
  invx g0132(.a(n432), .O(n433));
  orx  g0133(.a(n433), .b(n431), .O(n434));
  orx  g0134(.a(n434), .b(n421), .O(n435));
  invx g0135(.a(pi064), .O(n436));
  andx g0136(.a(n436), .b(pi079), .O(n437));
  andx g0137(.a(n437), .b(pi077), .O(n438));
  invx g0138(.a(n438), .O(n439));
  andx g0139(.a(n436), .b(n419), .O(n440));
  invx g0140(.a(n440), .O(n441));
  andx g0141(.a(pi007), .b(pi027), .O(n442));
  andx g0142(.a(pi005), .b(n312), .O(n443));
  orx  g0143(.a(n443), .b(pi026), .O(n444));
  orx  g0144(.a(n444), .b(n442), .O(n445));
  invx g0145(.a(pi034), .O(n446));
  andx g0146(.a(n446), .b(pi027), .O(n447));
  invx g0147(.a(pi003), .O(n448));
  andx g0148(.a(n448), .b(n312), .O(n449));
  orx  g0149(.a(n449), .b(n308), .O(n450));
  orx  g0150(.a(n450), .b(n447), .O(n451));
  andx g0151(.a(n451), .b(n445), .O(n452));
  orx  g0152(.a(n452), .b(n441), .O(n453));
  andx g0153(.a(n453), .b(n439), .O(n454));
  andx g0154(.a(n454), .b(n435), .O(po064));
  invx g0155(.a(po064), .O(n456));
  invx g0156(.a(pi119), .O(n457));
  andx g0157(.a(n457), .b(pi118), .O(n458));
  andx g0158(.a(n458), .b(n456), .O(n459));
  invx g0159(.a(pi040), .O(n460));
  invx g0160(.a(pi039), .O(po031));
  andx g0161(.a(po031), .b(pi061), .O(n462));
  invx g0162(.a(pi041), .O(n463));
  invx g0163(.a(pi061), .O(n464));
  andx g0164(.a(n464), .b(n463), .O(n465));
  orx  g0165(.a(n465), .b(n462), .O(n466));
  andx g0166(.a(n466), .b(n460), .O(n467));
  invx g0167(.a(n467), .O(n468));
  orx  g0168(.a(n466), .b(n460), .O(n469));
  andx g0169(.a(n469), .b(n468), .O(n470));
  invx g0170(.a(pi004), .O(n471));
  invx g0171(.a(pi038), .O(po014));
  andx g0172(.a(po014), .b(pi061), .O(n473));
  invx g0173(.a(pi045), .O(n474));
  andx g0174(.a(n474), .b(n464), .O(n475));
  orx  g0175(.a(n475), .b(n473), .O(n476));
  andx g0176(.a(n476), .b(n471), .O(n477));
  invx g0177(.a(n477), .O(n478));
  andx g0178(.a(n478), .b(n470), .O(n479));
  invx g0179(.a(n470), .O(n480));
  andx g0180(.a(n477), .b(n480), .O(n481));
  orx  g0181(.a(n481), .b(n421), .O(n482));
  orx  g0182(.a(n482), .b(n479), .O(n483));
  andx g0183(.a(n437), .b(pi076), .O(n484));
  invx g0184(.a(n484), .O(n485));
  andx g0185(.a(pi041), .b(pi007), .O(n486));
  andx g0186(.a(pi005), .b(n463), .O(n487));
  orx  g0187(.a(n487), .b(pi040), .O(n488));
  orx  g0188(.a(n488), .b(n486), .O(n489));
  andx g0189(.a(n446), .b(pi041), .O(n490));
  andx g0190(.a(n448), .b(n463), .O(n491));
  orx  g0191(.a(n491), .b(n460), .O(n492));
  orx  g0192(.a(n492), .b(n490), .O(n493));
  andx g0193(.a(n493), .b(n489), .O(n494));
  orx  g0194(.a(n494), .b(n441), .O(n495));
  andx g0195(.a(n495), .b(n485), .O(n496));
  andx g0196(.a(n496), .b(n483), .O(po025));
  invx g0197(.a(po025), .O(n498));
  invx g0198(.a(pi118), .O(n499));
  andx g0199(.a(n457), .b(n499), .O(n500));
  andx g0200(.a(n500), .b(n498), .O(n501));
  andx g0201(.a(pi119), .b(n499), .O(n502));
  andx g0202(.a(n502), .b(pi129), .O(n503));
  andx g0203(.a(pi119), .b(pi118), .O(n504));
  andx g0204(.a(n504), .b(pi128), .O(n505));
  orx  g0205(.a(n505), .b(n503), .O(n506));
  orx  g0206(.a(n506), .b(n501), .O(n507));
  orx  g0207(.a(n507), .b(n459), .O(n508));
  andx g0208(.a(n508), .b(pi120), .O(po002));
  invx g0209(.a(pi120), .O(n510));
  andx g0210(.a(n379), .b(n368), .O(n511));
  invx g0211(.a(n511), .O(n512));
  andx g0212(.a(n512), .b(n409), .O(n513));
  andx g0213(.a(n513), .b(n404), .O(n514));
  invx g0214(.a(n513), .O(n515));
  andx g0215(.a(n515), .b(n405), .O(n516));
  orx  g0216(.a(n516), .b(n514), .O(n517));
  andx g0217(.a(n375), .b(n367), .O(n518));
  invx g0218(.a(n518), .O(n519));
  andx g0219(.a(n519), .b(n410), .O(n520));
  invx g0220(.a(n520), .O(n521));
  invx g0221(.a(n394), .O(n522));
  andx g0222(.a(n413), .b(n522), .O(n523));
  orx  g0223(.a(n523), .b(n521), .O(n524));
  andx g0224(.a(n523), .b(n521), .O(n525));
  invx g0225(.a(n525), .O(n526));
  andx g0226(.a(n526), .b(n524), .O(n527));
  invx g0227(.a(n527), .O(n528));
  andx g0228(.a(n528), .b(n517), .O(n529));
  invx g0229(.a(n529), .O(n530));
  orx  g0230(.a(n528), .b(n517), .O(n531));
  andx g0231(.a(n531), .b(n530), .O(n532));
  orx  g0232(.a(n319), .b(pi026), .O(n533));
  andx g0233(.a(n533), .b(n315), .O(n534));
  andx g0234(.a(n427), .b(n534), .O(n535));
  andx g0235(.a(n342), .b(n340), .O(n536));
  invx g0236(.a(n332), .O(n537));
  andx g0237(.a(n537), .b(n307), .O(n538));
  andx g0238(.a(n538), .b(n536), .O(n539));
  andx g0239(.a(n539), .b(n535), .O(n540));
  orx  g0240(.a(n355), .b(n350), .O(n541));
  invx g0241(.a(n541), .O(n542));
  andx g0242(.a(n542), .b(n540), .O(n543));
  andx g0243(.a(n543), .b(pi033), .O(n544));
  orx  g0244(.a(n544), .b(n357), .O(n545));
  invx g0245(.a(n545), .O(n546));
  orx  g0246(.a(n546), .b(n532), .O(n547));
  andx g0247(.a(n411), .b(n391), .O(n548));
  invx g0248(.a(n548), .O(n549));
  andx g0249(.a(n549), .b(n412), .O(n550));
  andx g0250(.a(n550), .b(n404), .O(n551));
  invx g0251(.a(n551), .O(n552));
  orx  g0252(.a(n550), .b(n404), .O(n553));
  andx g0253(.a(n553), .b(n552), .O(n554));
  invx g0254(.a(n554), .O(n555));
  andx g0255(.a(n378), .b(n367), .O(n556));
  orx  g0256(.a(n556), .b(n511), .O(n557));
  andx g0257(.a(n557), .b(n555), .O(n558));
  invx g0258(.a(n558), .O(n559));
  orx  g0259(.a(n557), .b(n555), .O(n560));
  andx g0260(.a(n560), .b(n559), .O(n561));
  orx  g0261(.a(n561), .b(n545), .O(n562));
  andx g0262(.a(n562), .b(n547), .O(n563));
  invx g0263(.a(n563), .O(n564));
  orx  g0264(.a(n564), .b(n392), .O(n565));
  invx g0265(.a(n392), .O(n566));
  orx  g0266(.a(n563), .b(n566), .O(n567));
  andx g0267(.a(n567), .b(n565), .O(n568));
  invx g0268(.a(n568), .O(n569));
  orx  g0269(.a(pi022), .b(n311), .O(n570));
  andx g0270(.a(n304), .b(n570), .O(n571));
  andx g0271(.a(n571), .b(pi023), .O(n572));
  orx  g0272(.a(n320), .b(n572), .O(n573));
  andx g0273(.a(n537), .b(n329), .O(n574));
  andx g0274(.a(n574), .b(n573), .O(n575));
  andx g0275(.a(n333), .b(n424), .O(n576));
  orx  g0276(.a(n576), .b(n575), .O(n577));
  invx g0277(.a(n577), .O(n578));
  andx g0278(.a(n424), .b(n534), .O(n579));
  orx  g0279(.a(n579), .b(n573), .O(n580));
  andx g0280(.a(n537), .b(n580), .O(n581));
  orx  g0281(.a(n339), .b(n581), .O(n582));
  andx g0282(.a(n342), .b(n582), .O(n583));
  andx g0283(.a(n330), .b(n315), .O(n584));
  invx g0284(.a(n584), .O(n585));
  andx g0285(.a(n585), .b(n583), .O(n586));
  andx g0286(.a(n584), .b(n344), .O(n587));
  orx  g0287(.a(n587), .b(n586), .O(n588));
  andx g0288(.a(n588), .b(n578), .O(n589));
  orx  g0289(.a(n584), .b(n344), .O(n590));
  orx  g0290(.a(n585), .b(n583), .O(n591));
  andx g0291(.a(n591), .b(n590), .O(n592));
  andx g0292(.a(n592), .b(n577), .O(n593));
  orx  g0293(.a(n593), .b(n589), .O(n594));
  andx g0294(.a(n594), .b(n542), .O(n595));
  orx  g0295(.a(n592), .b(n577), .O(n596));
  orx  g0296(.a(n588), .b(n578), .O(n597));
  andx g0297(.a(n597), .b(n596), .O(n598));
  andx g0298(.a(n598), .b(n541), .O(n599));
  orx  g0299(.a(n599), .b(n595), .O(n600));
  andx g0300(.a(n426), .b(n322), .O(n601));
  orx  g0301(.a(n601), .b(n535), .O(n602));
  andx g0302(.a(n602), .b(n600), .O(n603));
  invx g0303(.a(n603), .O(n604));
  orx  g0304(.a(n602), .b(n600), .O(n605));
  andx g0305(.a(n605), .b(n604), .O(n606));
  orx  g0306(.a(n606), .b(pi033), .O(n607));
  invx g0307(.a(pi033), .O(n608));
  orx  g0308(.a(n594), .b(n427), .O(n609));
  invx g0309(.a(n535), .O(n610));
  orx  g0310(.a(n343), .b(n339), .O(n611));
  invx g0311(.a(n538), .O(n612));
  orx  g0312(.a(n612), .b(n611), .O(n613));
  orx  g0313(.a(n613), .b(n610), .O(n614));
  andx g0314(.a(n614), .b(n344), .O(n615));
  andx g0315(.a(n538), .b(n535), .O(n616));
  orx  g0316(.a(n616), .b(n581), .O(n617));
  andx g0317(.a(n617), .b(n615), .O(n618));
  orx  g0318(.a(n540), .b(n583), .O(n619));
  invx g0319(.a(n617), .O(n620));
  andx g0320(.a(n620), .b(n619), .O(n621));
  orx  g0321(.a(n621), .b(n618), .O(n622));
  andx g0322(.a(n584), .b(n610), .O(n623));
  orx  g0323(.a(n623), .b(n622), .O(n624));
  orx  g0324(.a(n620), .b(n619), .O(n625));
  orx  g0325(.a(n617), .b(n615), .O(n626));
  andx g0326(.a(n626), .b(n625), .O(n627));
  invx g0327(.a(n623), .O(n628));
  orx  g0328(.a(n628), .b(n627), .O(n629));
  andx g0329(.a(n629), .b(n624), .O(n630));
  orx  g0330(.a(n630), .b(n426), .O(n631));
  andx g0331(.a(n631), .b(n609), .O(n632));
  orx  g0332(.a(n632), .b(n322), .O(n633));
  andx g0333(.a(n598), .b(n426), .O(n634));
  andx g0334(.a(n628), .b(n627), .O(n635));
  andx g0335(.a(n623), .b(n622), .O(n636));
  orx  g0336(.a(n636), .b(n635), .O(n637));
  andx g0337(.a(n637), .b(n427), .O(n638));
  orx  g0338(.a(n638), .b(n634), .O(n639));
  orx  g0339(.a(n639), .b(n534), .O(n640));
  andx g0340(.a(n640), .b(n633), .O(n641));
  orx  g0341(.a(n641), .b(n542), .O(n642));
  andx g0342(.a(n639), .b(n534), .O(n643));
  andx g0343(.a(n632), .b(n322), .O(n644));
  orx  g0344(.a(n644), .b(n643), .O(n645));
  orx  g0345(.a(n645), .b(n541), .O(n646));
  andx g0346(.a(n646), .b(n642), .O(n647));
  orx  g0347(.a(n647), .b(n608), .O(n648));
  andx g0348(.a(n648), .b(n607), .O(n649));
  andx g0349(.a(n612), .b(n611), .O(n650));
  orx  g0350(.a(n650), .b(n539), .O(n651));
  andx g0351(.a(n651), .b(n649), .O(n652));
  invx g0352(.a(n607), .O(n653));
  andx g0353(.a(n645), .b(n541), .O(n654));
  andx g0354(.a(n641), .b(n542), .O(n655));
  orx  g0355(.a(n655), .b(n654), .O(n656));
  andx g0356(.a(n656), .b(pi033), .O(n657));
  orx  g0357(.a(n657), .b(n653), .O(n658));
  invx g0358(.a(n651), .O(n659));
  andx g0359(.a(n659), .b(n658), .O(n660));
  orx  g0360(.a(n660), .b(n652), .O(n661));
  orx  g0361(.a(n661), .b(n569), .O(n662));
  orx  g0362(.a(n659), .b(n658), .O(n663));
  orx  g0363(.a(n651), .b(n649), .O(n664));
  andx g0364(.a(n664), .b(n663), .O(n665));
  orx  g0365(.a(n665), .b(n568), .O(n666));
  andx g0366(.a(n666), .b(n420), .O(n667));
  andx g0367(.a(n667), .b(n662), .O(n668));
  invx g0368(.a(pi051), .O(n669));
  andx g0369(.a(n669), .b(pi024), .O(n670));
  invx g0370(.a(pi024), .O(n671));
  invx g0371(.a(pi050), .O(n672));
  andx g0372(.a(n672), .b(n671), .O(n673));
  orx  g0373(.a(n673), .b(pi023), .O(n674));
  orx  g0374(.a(n674), .b(n670), .O(n675));
  andx g0375(.a(pi046), .b(pi024), .O(n676));
  andx g0376(.a(pi047), .b(n671), .O(n677));
  orx  g0377(.a(n677), .b(n301), .O(n678));
  orx  g0378(.a(n678), .b(n676), .O(n679));
  andx g0379(.a(n679), .b(n675), .O(n680));
  andx g0380(.a(n669), .b(pi021), .O(n681));
  andx g0381(.a(n672), .b(n335), .O(n682));
  orx  g0382(.a(n682), .b(pi020), .O(n683));
  orx  g0383(.a(n683), .b(n681), .O(n684));
  andx g0384(.a(pi046), .b(pi021), .O(n685));
  invx g0385(.a(pi020), .O(n686));
  andx g0386(.a(pi047), .b(n335), .O(n687));
  orx  g0387(.a(n687), .b(n686), .O(n688));
  orx  g0388(.a(n688), .b(n685), .O(n689));
  andx g0389(.a(n689), .b(n684), .O(n690));
  invx g0390(.a(n690), .O(n691));
  andx g0391(.a(n669), .b(pi030), .O(n692));
  invx g0392(.a(pi030), .O(n693));
  andx g0393(.a(n672), .b(n693), .O(n694));
  orx  g0394(.a(n694), .b(pi031), .O(n695));
  orx  g0395(.a(n695), .b(n692), .O(n696));
  andx g0396(.a(pi046), .b(pi030), .O(n697));
  andx g0397(.a(pi047), .b(n693), .O(n698));
  orx  g0398(.a(n698), .b(n323), .O(n699));
  orx  g0399(.a(n699), .b(n697), .O(n700));
  andx g0400(.a(n700), .b(n696), .O(n701));
  andx g0401(.a(n701), .b(n691), .O(n702));
  invx g0402(.a(n702), .O(n703));
  orx  g0403(.a(n701), .b(n691), .O(n704));
  andx g0404(.a(n704), .b(n703), .O(n705));
  invx g0405(.a(n705), .O(n706));
  andx g0406(.a(n706), .b(n680), .O(n707));
  invx g0407(.a(n707), .O(n708));
  orx  g0408(.a(n706), .b(n680), .O(n709));
  andx g0409(.a(n709), .b(n708), .O(n710));
  invx g0410(.a(n710), .O(n711));
  andx g0411(.a(n669), .b(pi018), .O(n712));
  andx g0412(.a(n672), .b(n346), .O(n713));
  orx  g0413(.a(n713), .b(pi017), .O(n714));
  orx  g0414(.a(n714), .b(n712), .O(n715));
  andx g0415(.a(pi046), .b(pi018), .O(n716));
  andx g0416(.a(pi047), .b(n346), .O(n717));
  orx  g0417(.a(n717), .b(n353), .O(n718));
  orx  g0418(.a(n718), .b(n716), .O(n719));
  andx g0419(.a(n719), .b(n715), .O(n720));
  andx g0420(.a(n669), .b(pi027), .O(n721));
  andx g0421(.a(n672), .b(n312), .O(n722));
  orx  g0422(.a(n722), .b(pi026), .O(n723));
  orx  g0423(.a(n723), .b(n721), .O(n724));
  andx g0424(.a(pi046), .b(pi027), .O(n725));
  andx g0425(.a(pi047), .b(n312), .O(n726));
  orx  g0426(.a(n726), .b(n308), .O(n727));
  orx  g0427(.a(n727), .b(n725), .O(n728));
  andx g0428(.a(n728), .b(n724), .O(n729));
  invx g0429(.a(n729), .O(n730));
  andx g0430(.a(n730), .b(n720), .O(n731));
  invx g0431(.a(n731), .O(n732));
  orx  g0432(.a(n730), .b(n720), .O(n733));
  andx g0433(.a(n733), .b(n732), .O(n734));
  invx g0434(.a(n734), .O(n735));
  andx g0435(.a(n735), .b(n711), .O(n736));
  andx g0436(.a(n734), .b(n710), .O(n737));
  orx  g0437(.a(n737), .b(n736), .O(n738));
  invx g0438(.a(n738), .O(n739));
  andx g0439(.a(n669), .b(pi036), .O(n740));
  andx g0440(.a(n672), .b(n397), .O(n741));
  orx  g0441(.a(n741), .b(pi037), .O(n742));
  orx  g0442(.a(n742), .b(n740), .O(n743));
  andx g0443(.a(pi046), .b(pi036), .O(n744));
  andx g0444(.a(pi047), .b(n397), .O(n745));
  orx  g0445(.a(n745), .b(n395), .O(n746));
  orx  g0446(.a(n746), .b(n744), .O(n747));
  andx g0447(.a(n747), .b(n743), .O(n748));
  andx g0448(.a(n669), .b(pi009), .O(n749));
  andx g0449(.a(n672), .b(n359), .O(n750));
  orx  g0450(.a(n750), .b(pi010), .O(n751));
  orx  g0451(.a(n751), .b(n749), .O(n752));
  andx g0452(.a(pi046), .b(pi009), .O(n753));
  andx g0453(.a(pi047), .b(n359), .O(n754));
  orx  g0454(.a(n754), .b(n364), .O(n755));
  orx  g0455(.a(n755), .b(n753), .O(n756));
  andx g0456(.a(n756), .b(n752), .O(n757));
  invx g0457(.a(n757), .O(n758));
  andx g0458(.a(n758), .b(n748), .O(n759));
  invx g0459(.a(n748), .O(n760));
  andx g0460(.a(n757), .b(n760), .O(n761));
  orx  g0461(.a(n761), .b(n759), .O(n762));
  andx g0462(.a(n669), .b(pi015), .O(n763));
  andx g0463(.a(n672), .b(n383), .O(n764));
  orx  g0464(.a(n764), .b(pi014), .O(n765));
  orx  g0465(.a(n765), .b(n763), .O(n766));
  andx g0466(.a(pi046), .b(pi015), .O(n767));
  andx g0467(.a(pi047), .b(n383), .O(n768));
  orx  g0468(.a(n768), .b(n381), .O(n769));
  orx  g0469(.a(n769), .b(n767), .O(n770));
  andx g0470(.a(n770), .b(n766), .O(n771));
  andx g0471(.a(n669), .b(pi012), .O(n772));
  andx g0472(.a(n672), .b(n370), .O(n773));
  orx  g0473(.a(n773), .b(pi011), .O(n774));
  orx  g0474(.a(n774), .b(n772), .O(n775));
  andx g0475(.a(pi046), .b(pi012), .O(n776));
  andx g0476(.a(pi047), .b(n370), .O(n777));
  orx  g0477(.a(n777), .b(n376), .O(n778));
  orx  g0478(.a(n778), .b(n776), .O(n779));
  andx g0479(.a(n779), .b(n775), .O(n780));
  invx g0480(.a(n780), .O(n781));
  andx g0481(.a(n781), .b(n771), .O(n782));
  invx g0482(.a(n782), .O(n783));
  orx  g0483(.a(n781), .b(n771), .O(n784));
  andx g0484(.a(n784), .b(n783), .O(n785));
  invx g0485(.a(n785), .O(n786));
  andx g0486(.a(n786), .b(n762), .O(n787));
  invx g0487(.a(n787), .O(n788));
  orx  g0488(.a(n786), .b(n762), .O(n789));
  andx g0489(.a(n789), .b(n788), .O(n790));
  andx g0490(.a(n790), .b(n739), .O(n791));
  invx g0491(.a(n791), .O(n792));
  orx  g0492(.a(n790), .b(n739), .O(n793));
  andx g0493(.a(n793), .b(n440), .O(n794));
  andx g0494(.a(n794), .b(n792), .O(n795));
  orx  g0495(.a(n795), .b(pi079), .O(n796));
  orx  g0496(.a(n796), .b(n668), .O(n797));
  andx g0497(.a(pi091), .b(pi079), .O(n798));
  invx g0498(.a(n798), .O(n799));
  andx g0499(.a(n799), .b(n797), .O(n800));
  invx g0500(.a(pi121), .O(n801));
  andx g0501(.a(n801), .b(pi117), .O(n802));
  invx g0502(.a(n802), .O(n803));
  orx  g0503(.a(n803), .b(n800), .O(n804));
  invx g0504(.a(pi002), .O(n805));
  andx g0505(.a(n476), .b(n469), .O(n806));
  orx  g0506(.a(n806), .b(n467), .O(n807));
  invx g0507(.a(n807), .O(n808));
  invx g0508(.a(pi053), .O(n809));
  invx g0509(.a(pi054), .O(n810));
  andx g0510(.a(n810), .b(pi061), .O(n811));
  invx g0511(.a(pi052), .O(n812));
  andx g0512(.a(n812), .b(n464), .O(n813));
  orx  g0513(.a(n813), .b(n811), .O(n814));
  andx g0514(.a(n814), .b(n809), .O(n815));
  invx g0515(.a(n815), .O(n816));
  invx g0516(.a(n814), .O(n817));
  andx g0517(.a(n817), .b(pi053), .O(n818));
  invx g0518(.a(n818), .O(n819));
  andx g0519(.a(n819), .b(n816), .O(n820));
  invx g0520(.a(n820), .O(n821));
  andx g0521(.a(n821), .b(n808), .O(n822));
  andx g0522(.a(n820), .b(n807), .O(n823));
  orx  g0523(.a(n823), .b(n822), .O(n824));
  invx g0524(.a(n824), .O(n825));
  invx g0525(.a(pi044), .O(po105));
  andx g0526(.a(po105), .b(pi061), .O(n827));
  invx g0527(.a(pi042), .O(n828));
  andx g0528(.a(n828), .b(n464), .O(n829));
  orx  g0529(.a(n829), .b(n827), .O(n830));
  invx g0530(.a(n830), .O(n831));
  andx g0531(.a(n831), .b(pi043), .O(n832));
  invx g0532(.a(n832), .O(n833));
  andx g0533(.a(n833), .b(n807), .O(n834));
  invx g0534(.a(pi043), .O(n835));
  andx g0535(.a(n830), .b(n835), .O(n836));
  orx  g0536(.a(n836), .b(n834), .O(n837));
  andx g0537(.a(n837), .b(n470), .O(n838));
  invx g0538(.a(n837), .O(n839));
  andx g0539(.a(n839), .b(n480), .O(n840));
  orx  g0540(.a(n840), .b(n838), .O(n841));
  orx  g0541(.a(n841), .b(n825), .O(n842));
  andx g0542(.a(n841), .b(n825), .O(n843));
  invx g0543(.a(n843), .O(n844));
  andx g0544(.a(n844), .b(n842), .O(n845));
  invx g0545(.a(n845), .O(n846));
  invx g0546(.a(pi048), .O(n847));
  invx g0547(.a(pi049), .O(po015));
  andx g0548(.a(po015), .b(pi061), .O(n849));
  andx g0549(.a(n849), .b(n847), .O(n850));
  orx  g0550(.a(n850), .b(n837), .O(n851));
  invx g0551(.a(n849), .O(n852));
  andx g0552(.a(n852), .b(pi048), .O(n853));
  invx g0553(.a(n853), .O(n854));
  andx g0554(.a(n854), .b(n851), .O(n855));
  invx g0555(.a(n855), .O(n856));
  andx g0556(.a(n856), .b(n846), .O(n857));
  andx g0557(.a(n855), .b(n845), .O(n858));
  orx  g0558(.a(n858), .b(n857), .O(n859));
  andx g0559(.a(n859), .b(n805), .O(n860));
  invx g0560(.a(n860), .O(n861));
  andx g0561(.a(n806), .b(n468), .O(n862));
  invx g0562(.a(n836), .O(n863));
  andx g0563(.a(n863), .b(n833), .O(n864));
  orx  g0564(.a(n853), .b(n850), .O(n865));
  invx g0565(.a(n865), .O(n866));
  andx g0566(.a(n866), .b(n864), .O(n867));
  andx g0567(.a(n867), .b(n862), .O(n868));
  invx g0568(.a(n868), .O(n869));
  andx g0569(.a(n869), .b(n855), .O(n870));
  invx g0570(.a(n476), .O(n871));
  andx g0571(.a(n871), .b(n480), .O(n872));
  orx  g0572(.a(n872), .b(n862), .O(n873));
  andx g0573(.a(n873), .b(n870), .O(n874));
  orx  g0574(.a(n873), .b(n855), .O(n875));
  invx g0575(.a(n875), .O(n876));
  orx  g0576(.a(n876), .b(n874), .O(n877));
  andx g0577(.a(n863), .b(n468), .O(n878));
  andx g0578(.a(n833), .b(n467), .O(n879));
  orx  g0579(.a(n879), .b(n878), .O(n880));
  invx g0580(.a(n880), .O(n881));
  andx g0581(.a(n881), .b(n821), .O(n882));
  andx g0582(.a(n880), .b(n820), .O(n883));
  orx  g0583(.a(n883), .b(n882), .O(n884));
  orx  g0584(.a(n884), .b(n877), .O(n885));
  andx g0585(.a(n884), .b(n877), .O(n886));
  invx g0586(.a(n886), .O(n887));
  andx g0587(.a(n887), .b(n885), .O(n888));
  orx  g0588(.a(n888), .b(n805), .O(n889));
  andx g0589(.a(n889), .b(n861), .O(n890));
  andx g0590(.a(n856), .b(n816), .O(n891));
  orx  g0591(.a(n891), .b(n818), .O(n892));
  andx g0592(.a(n868), .b(n820), .O(n893));
  andx g0593(.a(n893), .b(pi002), .O(n894));
  orx  g0594(.a(n894), .b(n892), .O(n895));
  invx g0595(.a(n895), .O(n896));
  orx  g0596(.a(pi063), .b(n464), .O(n897));
  invx g0597(.a(pi059), .O(n898));
  andx g0598(.a(n898), .b(n464), .O(n899));
  invx g0599(.a(n899), .O(n900));
  andx g0600(.a(n900), .b(n897), .O(n901));
  andx g0601(.a(n901), .b(pi060), .O(n902));
  orx  g0602(.a(pi055), .b(n464), .O(n903));
  invx g0603(.a(pi057), .O(n904));
  andx g0604(.a(n904), .b(n464), .O(n905));
  invx g0605(.a(n905), .O(n906));
  andx g0606(.a(n906), .b(n903), .O(n907));
  andx g0607(.a(n907), .b(pi056), .O(n908));
  invx g0608(.a(pi060), .O(n909));
  invx g0609(.a(n901), .O(n910));
  andx g0610(.a(n910), .b(n909), .O(n911));
  orx  g0611(.a(n911), .b(n902), .O(n912));
  invx g0612(.a(n912), .O(n913));
  andx g0613(.a(n913), .b(n908), .O(n914));
  orx  g0614(.a(n914), .b(n902), .O(n915));
  orx  g0615(.a(pi062), .b(n464), .O(n916));
  invx g0616(.a(pi058), .O(n917));
  andx g0617(.a(n917), .b(n464), .O(n918));
  invx g0618(.a(n918), .O(n919));
  andx g0619(.a(n919), .b(n916), .O(n920));
  invx g0620(.a(n920), .O(n921));
  orx  g0621(.a(n921), .b(n915), .O(n922));
  invx g0622(.a(pi066), .O(po013));
  andx g0623(.a(po013), .b(pi061), .O(n924));
  invx g0624(.a(pi065), .O(n925));
  andx g0625(.a(n925), .b(n464), .O(n926));
  orx  g0626(.a(n926), .b(n924), .O(n927));
  invx g0627(.a(n927), .O(n928));
  orx  g0628(.a(n928), .b(n922), .O(n929));
  andx g0629(.a(n928), .b(n921), .O(n930));
  andx g0630(.a(n927), .b(n920), .O(n931));
  orx  g0631(.a(n931), .b(n930), .O(n932));
  invx g0632(.a(n932), .O(n933));
  andx g0633(.a(n933), .b(n922), .O(n934));
  invx g0634(.a(n934), .O(n935));
  andx g0635(.a(n935), .b(n929), .O(n936));
  invx g0636(.a(pi056), .O(n937));
  invx g0637(.a(n907), .O(n938));
  andx g0638(.a(n938), .b(n937), .O(n939));
  andx g0639(.a(n939), .b(n912), .O(n940));
  invx g0640(.a(n939), .O(n941));
  andx g0641(.a(n941), .b(n913), .O(n942));
  orx  g0642(.a(n942), .b(n940), .O(n943));
  andx g0643(.a(n943), .b(n936), .O(n944));
  invx g0644(.a(n944), .O(n945));
  orx  g0645(.a(n943), .b(n936), .O(n946));
  andx g0646(.a(n946), .b(n945), .O(n947));
  andx g0647(.a(n947), .b(n896), .O(n948));
  invx g0648(.a(n948), .O(n949));
  invx g0649(.a(n908), .O(n950));
  andx g0650(.a(n912), .b(n950), .O(n951));
  orx  g0651(.a(n951), .b(n914), .O(n952));
  orx  g0652(.a(n942), .b(n902), .O(n953));
  andx g0653(.a(n953), .b(n920), .O(n954));
  andx g0654(.a(n954), .b(n952), .O(n955));
  invx g0655(.a(n955), .O(n956));
  orx  g0656(.a(n954), .b(n952), .O(n957));
  andx g0657(.a(n957), .b(n956), .O(n958));
  invx g0658(.a(n958), .O(n959));
  andx g0659(.a(n959), .b(n928), .O(n960));
  andx g0660(.a(n958), .b(n927), .O(n961));
  orx  g0661(.a(n961), .b(n960), .O(n962));
  orx  g0662(.a(n962), .b(n896), .O(n963));
  andx g0663(.a(n963), .b(n949), .O(n964));
  invx g0664(.a(n964), .O(n965));
  andx g0665(.a(n965), .b(n890), .O(n966));
  invx g0666(.a(n890), .O(n967));
  andx g0667(.a(n964), .b(n967), .O(n968));
  orx  g0668(.a(n968), .b(n966), .O(n969));
  invx g0669(.a(n864), .O(n970));
  andx g0670(.a(n865), .b(n970), .O(n971));
  orx  g0671(.a(n971), .b(n867), .O(n972));
  andx g0672(.a(n972), .b(n969), .O(n973));
  invx g0673(.a(n973), .O(n974));
  orx  g0674(.a(n972), .b(n969), .O(n975));
  andx g0675(.a(n975), .b(n420), .O(n976));
  andx g0676(.a(n976), .b(n974), .O(n977));
  andx g0677(.a(n669), .b(pi059), .O(n978));
  andx g0678(.a(n672), .b(n898), .O(n979));
  orx  g0679(.a(n979), .b(pi060), .O(n980));
  orx  g0680(.a(n980), .b(n978), .O(n981));
  andx g0681(.a(pi046), .b(pi059), .O(n982));
  andx g0682(.a(pi047), .b(n898), .O(n983));
  orx  g0683(.a(n983), .b(n909), .O(n984));
  orx  g0684(.a(n984), .b(n982), .O(n985));
  andx g0685(.a(n985), .b(n981), .O(n986));
  invx g0686(.a(n986), .O(n987));
  andx g0687(.a(pi057), .b(n669), .O(n988));
  andx g0688(.a(n904), .b(n672), .O(n989));
  orx  g0689(.a(n989), .b(pi056), .O(n990));
  orx  g0690(.a(n990), .b(n988), .O(n991));
  andx g0691(.a(pi057), .b(pi046), .O(n992));
  andx g0692(.a(n904), .b(pi047), .O(n993));
  orx  g0693(.a(n993), .b(n937), .O(n994));
  orx  g0694(.a(n994), .b(n992), .O(n995));
  andx g0695(.a(n995), .b(n991), .O(n996));
  invx g0696(.a(n996), .O(n997));
  andx g0697(.a(n997), .b(n987), .O(n998));
  andx g0698(.a(n996), .b(n986), .O(n999));
  orx  g0699(.a(n999), .b(n998), .O(n1000));
  invx g0700(.a(n1000), .O(n1001));
  andx g0701(.a(n925), .b(n672), .O(n1002));
  andx g0702(.a(pi065), .b(n669), .O(n1003));
  orx  g0703(.a(n1003), .b(n1002), .O(n1004));
  invx g0704(.a(n1004), .O(n1005));
  invx g0705(.a(pi047), .O(n1006));
  andx g0706(.a(n917), .b(n1006), .O(n1007));
  invx g0707(.a(pi046), .O(n1008));
  andx g0708(.a(pi058), .b(n1008), .O(n1009));
  orx  g0709(.a(n1009), .b(n1007), .O(n1010));
  andx g0710(.a(n1010), .b(n1005), .O(n1011));
  invx g0711(.a(n1010), .O(n1012));
  andx g0712(.a(n1012), .b(n1004), .O(n1013));
  orx  g0713(.a(n1013), .b(n1011), .O(n1014));
  andx g0714(.a(n1014), .b(n1001), .O(n1015));
  invx g0715(.a(n1015), .O(n1016));
  orx  g0716(.a(n1014), .b(n1001), .O(n1017));
  andx g0717(.a(n1017), .b(n1016), .O(n1018));
  invx g0718(.a(n1018), .O(n1019));
  andx g0719(.a(pi042), .b(n669), .O(n1020));
  andx g0720(.a(n828), .b(n672), .O(n1021));
  orx  g0721(.a(n1021), .b(pi043), .O(n1022));
  orx  g0722(.a(n1022), .b(n1020), .O(n1023));
  andx g0723(.a(pi042), .b(pi046), .O(n1024));
  andx g0724(.a(n828), .b(pi047), .O(n1025));
  orx  g0725(.a(n1025), .b(n835), .O(n1026));
  orx  g0726(.a(n1026), .b(n1024), .O(n1027));
  andx g0727(.a(n1027), .b(n1023), .O(n1028));
  andx g0728(.a(n669), .b(pi041), .O(n1029));
  andx g0729(.a(n672), .b(n463), .O(n1030));
  orx  g0730(.a(n1030), .b(pi040), .O(n1031));
  orx  g0731(.a(n1031), .b(n1029), .O(n1032));
  andx g0732(.a(pi046), .b(pi041), .O(n1033));
  andx g0733(.a(pi047), .b(n463), .O(n1034));
  orx  g0734(.a(n1034), .b(n460), .O(n1035));
  orx  g0735(.a(n1035), .b(n1033), .O(n1036));
  andx g0736(.a(n1036), .b(n1032), .O(n1037));
  invx g0737(.a(n1037), .O(n1038));
  andx g0738(.a(n1038), .b(n1028), .O(n1039));
  invx g0739(.a(n1039), .O(n1040));
  orx  g0740(.a(n1038), .b(n1028), .O(n1041));
  andx g0741(.a(n1041), .b(n1040), .O(n1042));
  andx g0742(.a(pi052), .b(n669), .O(n1043));
  andx g0743(.a(n812), .b(n672), .O(n1044));
  orx  g0744(.a(n1044), .b(pi053), .O(n1045));
  orx  g0745(.a(n1045), .b(n1043), .O(n1046));
  andx g0746(.a(pi052), .b(pi046), .O(n1047));
  andx g0747(.a(n812), .b(pi047), .O(n1048));
  orx  g0748(.a(n1048), .b(n809), .O(n1049));
  orx  g0749(.a(n1049), .b(n1047), .O(n1050));
  andx g0750(.a(n1050), .b(n1046), .O(n1051));
  invx g0751(.a(n1051), .O(n1052));
  andx g0752(.a(n1006), .b(n474), .O(n1053));
  andx g0753(.a(n1008), .b(pi045), .O(n1054));
  orx  g0754(.a(n1054), .b(n1053), .O(n1055));
  invx g0755(.a(n1055), .O(n1056));
  andx g0756(.a(n1056), .b(n1052), .O(n1057));
  andx g0757(.a(n1055), .b(n1051), .O(n1058));
  orx  g0758(.a(n1058), .b(n1057), .O(n1059));
  andx g0759(.a(n1059), .b(n1042), .O(n1060));
  invx g0760(.a(n1060), .O(n1061));
  orx  g0761(.a(n1059), .b(n1042), .O(n1062));
  andx g0762(.a(n1062), .b(n1061), .O(n1063));
  invx g0763(.a(n1063), .O(n1064));
  andx g0764(.a(n847), .b(pi051), .O(n1065));
  andx g0765(.a(pi048), .b(n1008), .O(n1066));
  orx  g0766(.a(n1066), .b(n1065), .O(n1067));
  andx g0767(.a(n1067), .b(n1064), .O(n1068));
  invx g0768(.a(n1068), .O(n1069));
  orx  g0769(.a(n1067), .b(n1064), .O(n1070));
  andx g0770(.a(n1070), .b(n1069), .O(n1071));
  andx g0771(.a(n1071), .b(n1019), .O(n1072));
  invx g0772(.a(n1072), .O(n1073));
  orx  g0773(.a(n1071), .b(n1019), .O(n1074));
  andx g0774(.a(n1074), .b(n440), .O(n1075));
  andx g0775(.a(n1075), .b(n1073), .O(n1076));
  orx  g0776(.a(n1076), .b(pi079), .O(n1077));
  orx  g0777(.a(n1077), .b(n977), .O(n1078));
  andx g0778(.a(pi092), .b(pi079), .O(n1079));
  invx g0779(.a(n1079), .O(n1080));
  andx g0780(.a(n1080), .b(n1078), .O(n1081));
  invx g0781(.a(pi117), .O(n1082));
  andx g0782(.a(n801), .b(n1082), .O(n1083));
  invx g0783(.a(n1083), .O(n1084));
  orx  g0784(.a(n1084), .b(n1081), .O(n1085));
  invx g0785(.a(pi130), .O(n1086));
  andx g0786(.a(pi121), .b(n1082), .O(n1087));
  invx g0787(.a(n1087), .O(n1088));
  orx  g0788(.a(n1088), .b(n1086), .O(n1089));
  invx g0789(.a(pi131), .O(n1090));
  andx g0790(.a(pi121), .b(pi117), .O(n1091));
  invx g0791(.a(n1091), .O(n1092));
  orx  g0792(.a(n1092), .b(n1090), .O(n1093));
  andx g0793(.a(n1093), .b(n1089), .O(n1094));
  andx g0794(.a(n1094), .b(n1085), .O(n1095));
  andx g0795(.a(n1095), .b(n804), .O(n1096));
  orx  g0796(.a(n1096), .b(n510), .O(po003));
  andx g0797(.a(n432), .b(n315), .O(n1098));
  andx g0798(.a(n1098), .b(n612), .O(n1099));
  orx  g0799(.a(n1098), .b(n612), .O(n1100));
  invx g0800(.a(n1100), .O(n1101));
  orx  g0801(.a(n1101), .b(n1099), .O(n1102));
  orx  g0802(.a(n1102), .b(n421), .O(n1103));
  andx g0803(.a(n437), .b(pi078), .O(n1104));
  invx g0804(.a(n1104), .O(n1105));
  andx g0805(.a(pi007), .b(pi024), .O(n1106));
  andx g0806(.a(pi005), .b(n671), .O(n1107));
  orx  g0807(.a(n1107), .b(pi023), .O(n1108));
  orx  g0808(.a(n1108), .b(n1106), .O(n1109));
  andx g0809(.a(n446), .b(pi024), .O(n1110));
  andx g0810(.a(n448), .b(n671), .O(n1111));
  orx  g0811(.a(n1111), .b(n301), .O(n1112));
  orx  g0812(.a(n1112), .b(n1110), .O(n1113));
  andx g0813(.a(n1113), .b(n1109), .O(n1114));
  orx  g0814(.a(n1114), .b(n441), .O(n1115));
  andx g0815(.a(n1115), .b(n1105), .O(n1116));
  andx g0816(.a(n1116), .b(n1103), .O(po052));
  invx g0817(.a(po052), .O(n1118));
  andx g0818(.a(n1118), .b(n802), .O(n1119));
  andx g0819(.a(n871), .b(pi004), .O(n1120));
  invx g0820(.a(n1120), .O(n1121));
  andx g0821(.a(n1121), .b(n479), .O(n1122));
  invx g0822(.a(n1122), .O(n1123));
  andx g0823(.a(n1123), .b(n807), .O(n1124));
  andx g0824(.a(n1124), .b(n970), .O(n1125));
  invx g0825(.a(n1125), .O(n1126));
  orx  g0826(.a(n1124), .b(n970), .O(n1127));
  andx g0827(.a(n1127), .b(n420), .O(n1128));
  andx g0828(.a(n1128), .b(n1126), .O(n1129));
  invx g0829(.a(n1129), .O(n1130));
  andx g0830(.a(n437), .b(pi084), .O(n1131));
  invx g0831(.a(n1131), .O(n1132));
  andx g0832(.a(pi042), .b(pi007), .O(n1133));
  andx g0833(.a(n828), .b(pi005), .O(n1134));
  orx  g0834(.a(n1134), .b(pi043), .O(n1135));
  orx  g0835(.a(n1135), .b(n1133), .O(n1136));
  andx g0836(.a(pi042), .b(n446), .O(n1137));
  andx g0837(.a(n828), .b(n448), .O(n1138));
  orx  g0838(.a(n1138), .b(n835), .O(n1139));
  orx  g0839(.a(n1139), .b(n1137), .O(n1140));
  andx g0840(.a(n1140), .b(n1136), .O(n1141));
  orx  g0841(.a(n1141), .b(n441), .O(n1142));
  andx g0842(.a(n1142), .b(n1132), .O(n1143));
  andx g0843(.a(n1143), .b(n1130), .O(po043));
  invx g0844(.a(po043), .O(n1145));
  andx g0845(.a(n1145), .b(n1083), .O(n1146));
  andx g0846(.a(n1087), .b(pi132), .O(n1147));
  andx g0847(.a(n1091), .b(pi133), .O(n1148));
  orx  g0848(.a(n1148), .b(n1147), .O(n1149));
  orx  g0849(.a(n1149), .b(n1146), .O(n1150));
  orx  g0850(.a(n1150), .b(n1119), .O(n1151));
  andx g0851(.a(n1151), .b(pi120), .O(po004));
  invx g0852(.a(n915), .O(n1153));
  andx g0853(.a(n934), .b(n1153), .O(n1154));
  invx g0854(.a(n1154), .O(n1155));
  andx g0855(.a(n942), .b(n950), .O(n1156));
  andx g0856(.a(n1156), .b(n1154), .O(n1157));
  andx g0857(.a(n1157), .b(n892), .O(n1158));
  orx  g0858(.a(n1158), .b(n1155), .O(po005));
  andx g0859(.a(n543), .b(n406), .O(po006));
  andx g0860(.a(n1157), .b(n893), .O(po007));
  andx g0861(.a(n1100), .b(n307), .O(n1162));
  andx g0862(.a(n1162), .b(n536), .O(n1163));
  invx g0863(.a(n1163), .O(n1164));
  andx g0864(.a(n1164), .b(n619), .O(n1165));
  andx g0865(.a(n1165), .b(n542), .O(n1166));
  invx g0866(.a(n1166), .O(n1167));
  andx g0867(.a(n1167), .b(n351), .O(n1168));
  andx g0868(.a(n1168), .b(n413), .O(n1169));
  orx  g0869(.a(n1169), .b(n523), .O(n1170));
  invx g0870(.a(n1170), .O(n1171));
  andx g0871(.a(n1171), .b(n404), .O(n1172));
  andx g0872(.a(n1170), .b(n405), .O(n1173));
  orx  g0873(.a(n1173), .b(n1172), .O(n1174));
  andx g0874(.a(n1174), .b(n420), .O(n1175));
  andx g0875(.a(n437), .b(pi083), .O(n1176));
  andx g0876(.a(n760), .b(n440), .O(n1177));
  orx  g0877(.a(n1177), .b(n1176), .O(n1178));
  orx  g0878(.a(n1178), .b(n1175), .O(n1179));
  andx g0879(.a(n1179), .b(n802), .O(n1180));
  andx g0880(.a(n1122), .b(n864), .O(n1181));
  orx  g0881(.a(n1181), .b(n839), .O(n1182));
  invx g0882(.a(n1182), .O(n1183));
  andx g0883(.a(n1183), .b(n866), .O(n1184));
  orx  g0884(.a(n1184), .b(n870), .O(n1185));
  invx g0885(.a(n1185), .O(n1186));
  andx g0886(.a(n1186), .b(n820), .O(n1187));
  invx g0887(.a(n1187), .O(n1188));
  andx g0888(.a(n1188), .b(n819), .O(n1189));
  andx g0889(.a(n1189), .b(n1153), .O(n1190));
  invx g0890(.a(n1190), .O(n1191));
  andx g0891(.a(n1191), .b(n953), .O(n1192));
  andx g0892(.a(n1192), .b(n927), .O(n1193));
  invx g0893(.a(n1193), .O(n1194));
  orx  g0894(.a(n1192), .b(n933), .O(n1195));
  andx g0895(.a(n1195), .b(n1194), .O(n1196));
  andx g0896(.a(n1196), .b(n420), .O(n1197));
  andx g0897(.a(n437), .b(pi072), .O(n1198));
  andx g0898(.a(n1005), .b(n440), .O(n1199));
  orx  g0899(.a(n1199), .b(n1198), .O(n1200));
  orx  g0900(.a(n1200), .b(n1197), .O(n1201));
  andx g0901(.a(n1201), .b(n1083), .O(n1202));
  andx g0902(.a(n1087), .b(pi134), .O(n1203));
  andx g0903(.a(n1091), .b(pi135), .O(n1204));
  orx  g0904(.a(n1204), .b(n1203), .O(n1205));
  orx  g0905(.a(n1205), .b(n1202), .O(n1206));
  orx  g0906(.a(n1206), .b(n1180), .O(n1207));
  andx g0907(.a(n1207), .b(pi120), .O(po008));
  invx g0908(.a(pi158), .O(n1209));
  andx g0909(.a(n1209), .b(pi159), .O(n1210));
  invx g0910(.a(pi159), .O(n1211));
  invx g0911(.a(pi157), .O(n1212));
  andx g0912(.a(n1212), .b(n1211), .O(n1213));
  invx g0913(.a(pi155), .O(n1214));
  invx g0914(.a(pi154), .O(n1215));
  orx  g0915(.a(n1215), .b(n1214), .O(po071));
  orx  g0916(.a(po071), .b(n1213), .O(n1217));
  orx  g0917(.a(n1217), .b(n1210), .O(po009));
  andx g0918(.a(n1196), .b(pi071), .O(n1219));
  invx g0919(.a(pi070), .O(n1220));
  invx g0920(.a(pi071), .O(n1221));
  andx g0921(.a(n1221), .b(pi072), .O(n1222));
  orx  g0922(.a(n1222), .b(n1220), .O(n1223));
  orx  g0923(.a(n1223), .b(n1219), .O(n1224));
  andx g0924(.a(n928), .b(pi069), .O(n1225));
  invx g0925(.a(pi069), .O(n1226));
  andx g0926(.a(n927), .b(n1226), .O(n1227));
  orx  g0927(.a(n1227), .b(n1225), .O(n1228));
  andx g0928(.a(n1228), .b(pi071), .O(n1229));
  andx g0929(.a(n1005), .b(n1221), .O(n1230));
  orx  g0930(.a(n1230), .b(pi070), .O(n1231));
  orx  g0931(.a(n1231), .b(n1229), .O(n1232));
  invx g0932(.a(pi145), .O(n1233));
  invx g0933(.a(pi144), .O(n1234));
  orx  g0934(.a(n1234), .b(n1233), .O(n1235));
  andx g0935(.a(n1235), .b(n1232), .O(n1236));
  andx g0936(.a(n1236), .b(n1224), .O(po010));
  invx g0937(.a(n380), .O(n1238));
  andx g0938(.a(n1168), .b(n1238), .O(n1239));
  invx g0939(.a(n1168), .O(n1240));
  andx g0940(.a(n1240), .b(n380), .O(n1241));
  orx  g0941(.a(n1241), .b(n1239), .O(n1242));
  orx  g0942(.a(n1242), .b(n421), .O(n1243));
  andx g0943(.a(n437), .b(pi073), .O(n1244));
  invx g0944(.a(n1244), .O(n1245));
  andx g0945(.a(pi007), .b(pi012), .O(n1246));
  andx g0946(.a(pi005), .b(n370), .O(n1247));
  orx  g0947(.a(n1247), .b(pi011), .O(n1248));
  orx  g0948(.a(n1248), .b(n1246), .O(n1249));
  andx g0949(.a(n446), .b(pi012), .O(n1250));
  andx g0950(.a(n448), .b(n370), .O(n1251));
  orx  g0951(.a(n1251), .b(n376), .O(n1252));
  orx  g0952(.a(n1252), .b(n1250), .O(n1253));
  andx g0953(.a(n1253), .b(n1249), .O(n1254));
  orx  g0954(.a(n1254), .b(n441), .O(n1255));
  andx g0955(.a(n1255), .b(n1245), .O(n1256));
  andx g0956(.a(n1256), .b(n1243), .O(po011));
  orx  g0957(.a(n1241), .b(n374), .O(n1258));
  orx  g0958(.a(n1258), .b(n368), .O(n1259));
  andx g0959(.a(n1258), .b(n368), .O(n1260));
  invx g0960(.a(n1260), .O(n1261));
  andx g0961(.a(n1261), .b(n1259), .O(n1262));
  andx g0962(.a(n1262), .b(n420), .O(n1263));
  andx g0963(.a(n437), .b(pi075), .O(n1264));
  invx g0964(.a(n1264), .O(n1265));
  andx g0965(.a(pi007), .b(pi009), .O(n1266));
  andx g0966(.a(pi005), .b(n359), .O(n1267));
  orx  g0967(.a(n1267), .b(pi010), .O(n1268));
  orx  g0968(.a(n1268), .b(n1266), .O(n1269));
  andx g0969(.a(n446), .b(pi009), .O(n1270));
  andx g0970(.a(n448), .b(n359), .O(n1271));
  orx  g0971(.a(n1271), .b(n364), .O(n1272));
  orx  g0972(.a(n1272), .b(n1270), .O(n1273));
  andx g0973(.a(n1273), .b(n1269), .O(n1274));
  orx  g0974(.a(n1274), .b(n441), .O(n1275));
  andx g0975(.a(n1275), .b(n1265), .O(n1276));
  invx g0976(.a(n1276), .O(n1277));
  orx  g0977(.a(n1277), .b(n1263), .O(n1278));
  andx g0978(.a(n1278), .b(n458), .O(n1279));
  invx g0979(.a(n1189), .O(n1280));
  andx g0980(.a(n1280), .b(n943), .O(n1281));
  andx g0981(.a(n1189), .b(n952), .O(n1282));
  orx  g0982(.a(n1282), .b(n1281), .O(n1283));
  orx  g0983(.a(n1283), .b(n421), .O(n1284));
  andx g0984(.a(n437), .b(pi074), .O(n1285));
  andx g0985(.a(n987), .b(n440), .O(n1286));
  orx  g0986(.a(n1286), .b(n1285), .O(n1287));
  invx g0987(.a(n1287), .O(n1288));
  andx g0988(.a(n1288), .b(n1284), .O(po120));
  invx g0989(.a(po120), .O(n1290));
  andx g0990(.a(n1290), .b(n500), .O(n1291));
  andx g0991(.a(n502), .b(pi126), .O(n1292));
  andx g0992(.a(n504), .b(pi127), .O(n1293));
  orx  g0993(.a(n1293), .b(n1292), .O(n1294));
  orx  g0994(.a(n1294), .b(n1291), .O(n1295));
  orx  g0995(.a(n1295), .b(n1279), .O(n1296));
  andx g0996(.a(n1296), .b(pi120), .O(po016));
  andx g0997(.a(n1121), .b(n478), .O(n1298));
  orx  g0998(.a(n1298), .b(n421), .O(n1299));
  andx g0999(.a(n437), .b(pi081), .O(n1300));
  andx g1000(.a(n1055), .b(n440), .O(n1301));
  orx  g1001(.a(n1301), .b(n1300), .O(n1302));
  invx g1002(.a(n1302), .O(n1303));
  andx g1003(.a(n1303), .b(n1299), .O(po017));
  invx g1004(.a(pi125), .O(n1305));
  andx g1005(.a(pi124), .b(n1305), .O(n1306));
  andx g1006(.a(n1306), .b(n1118), .O(n1307));
  invx g1007(.a(pi124), .O(n1308));
  andx g1008(.a(n1308), .b(n1305), .O(n1309));
  andx g1009(.a(n1309), .b(n1145), .O(n1310));
  andx g1010(.a(n1308), .b(pi125), .O(n1311));
  andx g1011(.a(n1311), .b(pi095), .O(n1312));
  andx g1012(.a(pi124), .b(pi125), .O(n1313));
  andx g1013(.a(n1313), .b(pi101), .O(n1314));
  orx  g1014(.a(n1314), .b(n1312), .O(n1315));
  orx  g1015(.a(n1315), .b(n1310), .O(n1316));
  orx  g1016(.a(n1316), .b(n1307), .O(po018));
  orx  g1017(.a(n427), .b(pi032), .O(n1318));
  andx g1018(.a(n1318), .b(n429), .O(n1319));
  andx g1019(.a(n1319), .b(n420), .O(n1320));
  invx g1020(.a(n1320), .O(n1321));
  andx g1021(.a(n437), .b(pi080), .O(n1322));
  invx g1022(.a(n1322), .O(n1323));
  andx g1023(.a(pi007), .b(pi030), .O(n1324));
  andx g1024(.a(pi005), .b(n693), .O(n1325));
  orx  g1025(.a(n1325), .b(pi031), .O(n1326));
  orx  g1026(.a(n1326), .b(n1324), .O(n1327));
  andx g1027(.a(n446), .b(pi030), .O(n1328));
  andx g1028(.a(n448), .b(n693), .O(n1329));
  orx  g1029(.a(n1329), .b(n323), .O(n1330));
  orx  g1030(.a(n1330), .b(n1328), .O(n1331));
  andx g1031(.a(n1331), .b(n1327), .O(n1332));
  orx  g1032(.a(n1332), .b(n441), .O(n1333));
  andx g1033(.a(n1333), .b(n1323), .O(n1334));
  andx g1034(.a(n1334), .b(n1321), .O(po051));
  invx g1035(.a(po051), .O(n1336));
  andx g1036(.a(n1336), .b(n1306), .O(n1337));
  invx g1037(.a(po017), .O(n1338));
  andx g1038(.a(n1309), .b(n1338), .O(n1339));
  andx g1039(.a(n1311), .b(pi110), .O(n1340));
  andx g1040(.a(n1313), .b(pi102), .O(n1341));
  orx  g1041(.a(n1341), .b(n1340), .O(n1342));
  orx  g1042(.a(n1342), .b(n1339), .O(n1343));
  orx  g1043(.a(n1343), .b(n1337), .O(po019));
  invx g1044(.a(pi122), .O(n1345));
  andx g1045(.a(n1345), .b(pi123), .O(n1346));
  andx g1046(.a(n1346), .b(n456), .O(n1347));
  invx g1047(.a(pi123), .O(n1348));
  andx g1048(.a(n1345), .b(n1348), .O(n1349));
  andx g1049(.a(n1349), .b(n498), .O(n1350));
  andx g1050(.a(pi122), .b(n1348), .O(n1351));
  andx g1051(.a(n1351), .b(pi096), .O(n1352));
  andx g1052(.a(pi122), .b(pi123), .O(n1353));
  andx g1053(.a(n1353), .b(pi097), .O(n1354));
  orx  g1054(.a(n1354), .b(n1352), .O(n1355));
  orx  g1055(.a(n1355), .b(n1350), .O(n1356));
  orx  g1056(.a(n1356), .b(n1347), .O(po020));
  andx g1057(.a(n400), .b(n377), .O(n1358));
  andx g1058(.a(n401), .b(n373), .O(n1359));
  orx  g1059(.a(n1359), .b(n1358), .O(n1360));
  invx g1060(.a(n1360), .O(n1361));
  andx g1061(.a(pi001), .b(pi028), .O(n1362));
  andx g1062(.a(pi006), .b(n311), .O(n1363));
  orx  g1063(.a(n1363), .b(n1362), .O(n1364));
  invx g1064(.a(n1364), .O(n1365));
  andx g1065(.a(n1365), .b(n365), .O(n1366));
  andx g1066(.a(n1364), .b(n362), .O(n1367));
  orx  g1067(.a(n1367), .b(n1366), .O(n1368));
  andx g1068(.a(n1368), .b(n387), .O(n1369));
  invx g1069(.a(n1369), .O(n1370));
  orx  g1070(.a(n1368), .b(n387), .O(n1371));
  andx g1071(.a(n1371), .b(n1370), .O(n1372));
  invx g1072(.a(n1372), .O(n1373));
  andx g1073(.a(n1373), .b(n1361), .O(n1374));
  andx g1074(.a(n1372), .b(n1360), .O(n1375));
  orx  g1075(.a(n1375), .b(n1374), .O(n1376));
  andx g1076(.a(n314), .b(n571), .O(n1377));
  andx g1077(.a(n319), .b(n306), .O(n1378));
  orx  g1078(.a(n1378), .b(n1377), .O(n1379));
  invx g1079(.a(n338), .O(n1380));
  andx g1080(.a(n1380), .b(n423), .O(n1381));
  andx g1081(.a(n338), .b(n328), .O(n1382));
  orx  g1082(.a(n1382), .b(n1381), .O(n1383));
  andx g1083(.a(n1383), .b(n1379), .O(n1384));
  invx g1084(.a(n1384), .O(n1385));
  orx  g1085(.a(n1383), .b(n1379), .O(n1386));
  andx g1086(.a(n1386), .b(n1385), .O(n1387));
  andx g1087(.a(n1387), .b(n354), .O(n1388));
  invx g1088(.a(n1388), .O(n1389));
  orx  g1089(.a(n1387), .b(n354), .O(n1390));
  andx g1090(.a(n1390), .b(n1389), .O(n1391));
  invx g1091(.a(n1391), .O(n1392));
  andx g1092(.a(n1392), .b(n1376), .O(n1393));
  invx g1093(.a(n1393), .O(n1394));
  orx  g1094(.a(n1392), .b(n1376), .O(n1395));
  andx g1095(.a(n1395), .b(n1394), .O(n1396));
  invx g1096(.a(n1396), .O(po021));
  invx g1097(.a(pi176), .O(po022));
  andx g1098(.a(n1278), .b(n802), .O(n1399));
  andx g1099(.a(n1290), .b(n1083), .O(n1400));
  andx g1100(.a(n1087), .b(pi126), .O(n1401));
  andx g1101(.a(n1091), .b(pi127), .O(n1402));
  orx  g1102(.a(n1402), .b(n1401), .O(n1403));
  orx  g1103(.a(n1403), .b(n1400), .O(n1404));
  orx  g1104(.a(n1404), .b(n1399), .O(n1405));
  andx g1105(.a(n1405), .b(pi120), .O(po023));
  orx  g1106(.a(n1162), .b(n536), .O(n1407));
  andx g1107(.a(n1407), .b(n1164), .O(n1408));
  orx  g1108(.a(n1408), .b(n421), .O(n1409));
  andx g1109(.a(n437), .b(pi082), .O(n1410));
  invx g1110(.a(n1410), .O(n1411));
  andx g1111(.a(pi007), .b(pi021), .O(n1412));
  andx g1112(.a(pi005), .b(n335), .O(n1413));
  orx  g1113(.a(n1413), .b(pi020), .O(n1414));
  orx  g1114(.a(n1414), .b(n1412), .O(n1415));
  andx g1115(.a(n446), .b(pi021), .O(n1416));
  andx g1116(.a(n448), .b(n335), .O(n1417));
  orx  g1117(.a(n1417), .b(n686), .O(n1418));
  orx  g1118(.a(n1418), .b(n1416), .O(n1419));
  andx g1119(.a(n1419), .b(n1415), .O(n1420));
  orx  g1120(.a(n1420), .b(n441), .O(n1421));
  andx g1121(.a(n1421), .b(n1411), .O(n1422));
  andx g1122(.a(n1422), .b(n1409), .O(po103));
  invx g1123(.a(po103), .O(n1424));
  andx g1124(.a(n1424), .b(n1346), .O(n1425));
  andx g1125(.a(n1182), .b(n865), .O(n1426));
  orx  g1126(.a(n1426), .b(n1184), .O(n1427));
  andx g1127(.a(n1427), .b(n420), .O(n1428));
  andx g1128(.a(n437), .b(pi087), .O(n1429));
  invx g1129(.a(pi007), .O(n1430));
  andx g1130(.a(n847), .b(n1430), .O(n1431));
  andx g1131(.a(pi048), .b(pi034), .O(n1432));
  orx  g1132(.a(n1432), .b(n1431), .O(n1433));
  andx g1133(.a(n1433), .b(n440), .O(n1434));
  orx  g1134(.a(n1434), .b(n1429), .O(n1435));
  orx  g1135(.a(n1435), .b(n1428), .O(n1436));
  andx g1136(.a(n1436), .b(n1349), .O(n1437));
  andx g1137(.a(n1351), .b(pi113), .O(n1438));
  andx g1138(.a(n1353), .b(pi114), .O(n1439));
  orx  g1139(.a(n1439), .b(n1438), .O(n1440));
  orx  g1140(.a(n1440), .b(n1437), .O(n1441));
  orx  g1141(.a(n1441), .b(n1425), .O(po024));
  andx g1142(.a(n1168), .b(n411), .O(n1443));
  orx  g1143(.a(n1443), .b(n513), .O(n1444));
  invx g1144(.a(n1444), .O(n1445));
  andx g1145(.a(n1445), .b(n566), .O(n1446));
  andx g1146(.a(n1444), .b(n392), .O(n1447));
  orx  g1147(.a(n1447), .b(n1446), .O(n1448));
  andx g1148(.a(n1448), .b(n420), .O(n1449));
  andx g1149(.a(n437), .b(pi088), .O(n1450));
  invx g1150(.a(n1450), .O(n1451));
  andx g1151(.a(pi007), .b(pi015), .O(n1452));
  andx g1152(.a(pi005), .b(n383), .O(n1453));
  orx  g1153(.a(n1453), .b(pi014), .O(n1454));
  orx  g1154(.a(n1454), .b(n1452), .O(n1455));
  andx g1155(.a(n446), .b(pi015), .O(n1456));
  andx g1156(.a(n448), .b(n383), .O(n1457));
  orx  g1157(.a(n1457), .b(n381), .O(n1458));
  orx  g1158(.a(n1458), .b(n1456), .O(n1459));
  andx g1159(.a(n1459), .b(n1455), .O(n1460));
  orx  g1160(.a(n1460), .b(n441), .O(n1461));
  andx g1161(.a(n1461), .b(n1451), .O(n1462));
  invx g1162(.a(n1462), .O(n1463));
  orx  g1163(.a(n1463), .b(n1449), .O(n1464));
  andx g1164(.a(n1464), .b(n1346), .O(n1465));
  andx g1165(.a(n1191), .b(n954), .O(n1466));
  orx  g1166(.a(n1192), .b(n920), .O(n1467));
  invx g1167(.a(n1467), .O(n1468));
  orx  g1168(.a(n1468), .b(n1466), .O(n1469));
  andx g1169(.a(n1469), .b(n420), .O(n1470));
  andx g1170(.a(n437), .b(pi085), .O(n1471));
  andx g1171(.a(n1010), .b(n440), .O(n1472));
  orx  g1172(.a(n1472), .b(n1471), .O(n1473));
  orx  g1173(.a(n1473), .b(n1470), .O(n1474));
  andx g1174(.a(n1474), .b(n1349), .O(n1475));
  andx g1175(.a(n1351), .b(pi098), .O(n1476));
  andx g1176(.a(n1353), .b(pi109), .O(n1477));
  orx  g1177(.a(n1477), .b(n1476), .O(n1478));
  orx  g1178(.a(n1478), .b(n1475), .O(n1479));
  orx  g1179(.a(n1479), .b(n1465), .O(po032));
  andx g1180(.a(n1346), .b(n1118), .O(n1481));
  andx g1181(.a(n1349), .b(n1145), .O(n1482));
  andx g1182(.a(n1351), .b(pi095), .O(n1483));
  andx g1183(.a(n1353), .b(pi101), .O(n1484));
  orx  g1184(.a(n1484), .b(n1483), .O(n1485));
  orx  g1185(.a(n1485), .b(n1482), .O(n1486));
  orx  g1186(.a(n1486), .b(n1481), .O(po033));
  andx g1187(.a(n1336), .b(n458), .O(n1488));
  andx g1188(.a(n1338), .b(n500), .O(n1489));
  andx g1189(.a(n502), .b(pi136), .O(n1490));
  andx g1190(.a(n504), .b(pi137), .O(n1491));
  orx  g1191(.a(n1491), .b(n1490), .O(n1492));
  orx  g1192(.a(n1492), .b(n1489), .O(n1493));
  orx  g1193(.a(n1493), .b(n1488), .O(n1494));
  andx g1194(.a(n1494), .b(pi120), .O(po034));
  andx g1195(.a(n1306), .b(n1179), .O(n1496));
  andx g1196(.a(n1309), .b(n1201), .O(n1497));
  andx g1197(.a(n1311), .b(pi104), .O(n1498));
  andx g1198(.a(n1313), .b(pi108), .O(n1499));
  orx  g1199(.a(n1499), .b(n1498), .O(n1500));
  orx  g1200(.a(n1500), .b(n1497), .O(n1501));
  orx  g1201(.a(n1501), .b(n1496), .O(po035));
  invx g1202(.a(pi170), .O(po036));
  andx g1203(.a(pi052), .b(pi007), .O(n1504));
  andx g1204(.a(n812), .b(pi005), .O(n1505));
  orx  g1205(.a(n1505), .b(pi053), .O(n1506));
  orx  g1206(.a(n1506), .b(n1504), .O(n1507));
  andx g1207(.a(pi052), .b(n446), .O(n1508));
  andx g1208(.a(n812), .b(n448), .O(n1509));
  orx  g1209(.a(n1509), .b(n809), .O(n1510));
  orx  g1210(.a(n1510), .b(n1508), .O(n1511));
  andx g1211(.a(n1511), .b(n1507), .O(n1512));
  invx g1212(.a(n1433), .O(n1513));
  andx g1213(.a(n1513), .b(n1056), .O(n1514));
  andx g1214(.a(n1514), .b(n1013), .O(n1515));
  andx g1215(.a(n1515), .b(n1512), .O(n1516));
  andx g1216(.a(n1141), .b(n494), .O(n1517));
  andx g1217(.a(n1517), .b(n1516), .O(n1518));
  andx g1218(.a(n1518), .b(n999), .O(po038));
  andx g1219(.a(pi147), .b(pi146), .O(po039));
  invx g1220(.a(pi153), .O(n1521));
  andx g1221(.a(n1521), .b(pi159), .O(n1522));
  invx g1222(.a(pi152), .O(n1523));
  andx g1223(.a(n1523), .b(n1211), .O(n1524));
  orx  g1224(.a(n1524), .b(n1522), .O(n1525));
  orx  g1225(.a(n1525), .b(po071), .O(po040));
  invx g1226(.a(po011), .O(n1527));
  andx g1227(.a(n1306), .b(n1527), .O(n1528));
  andx g1228(.a(n941), .b(n950), .O(n1529));
  invx g1229(.a(n1529), .O(n1530));
  andx g1230(.a(n1530), .b(n1189), .O(n1531));
  andx g1231(.a(n1529), .b(n1280), .O(n1532));
  orx  g1232(.a(n1532), .b(n1531), .O(n1533));
  orx  g1233(.a(n1533), .b(n421), .O(n1534));
  andx g1234(.a(n437), .b(pi090), .O(n1535));
  andx g1235(.a(n997), .b(n440), .O(n1536));
  orx  g1236(.a(n1536), .b(n1535), .O(n1537));
  invx g1237(.a(n1537), .O(n1538));
  andx g1238(.a(n1538), .b(n1534), .O(po081));
  invx g1239(.a(po081), .O(n1540));
  andx g1240(.a(n1540), .b(n1309), .O(n1541));
  andx g1241(.a(n1311), .b(pi107), .O(n1542));
  andx g1242(.a(n1313), .b(pi106), .O(n1543));
  orx  g1243(.a(n1543), .b(n1542), .O(n1544));
  orx  g1244(.a(n1544), .b(n1541), .O(n1545));
  orx  g1245(.a(n1545), .b(n1528), .O(po041));
  invx g1246(.a(n662), .O(n1547));
  andx g1247(.a(n661), .b(n569), .O(n1548));
  orx  g1248(.a(n1548), .b(n421), .O(n1549));
  orx  g1249(.a(n1549), .b(n1547), .O(n1550));
  invx g1250(.a(n796), .O(n1551));
  andx g1251(.a(n1551), .b(n1550), .O(n1552));
  orx  g1252(.a(n798), .b(n1552), .O(n1553));
  andx g1253(.a(n1306), .b(n1553), .O(n1554));
  invx g1254(.a(n1081), .O(n1555));
  andx g1255(.a(n1309), .b(n1555), .O(n1556));
  andx g1256(.a(n1311), .b(pi105), .O(n1557));
  andx g1257(.a(n1313), .b(pi103), .O(n1558));
  orx  g1258(.a(n1558), .b(n1557), .O(n1559));
  orx  g1259(.a(n1559), .b(n1556), .O(n1560));
  orx  g1260(.a(n1560), .b(n1554), .O(po042));
  andx g1261(.a(n1336), .b(n802), .O(n1562));
  andx g1262(.a(n1338), .b(n1083), .O(n1563));
  andx g1263(.a(n1087), .b(pi136), .O(n1564));
  andx g1264(.a(n1091), .b(pi137), .O(n1565));
  orx  g1265(.a(n1565), .b(n1564), .O(n1566));
  orx  g1266(.a(n1566), .b(n1563), .O(n1567));
  orx  g1267(.a(n1567), .b(n1562), .O(n1568));
  andx g1268(.a(n1568), .b(pi120), .O(po044));
  andx g1269(.a(n1424), .b(n802), .O(n1570));
  andx g1270(.a(n1436), .b(n1083), .O(n1571));
  andx g1271(.a(n1087), .b(pi116), .O(n1572));
  andx g1272(.a(n1091), .b(pi115), .O(n1573));
  orx  g1273(.a(n1573), .b(n1572), .O(n1574));
  orx  g1274(.a(n1574), .b(n1571), .O(n1575));
  orx  g1275(.a(n1575), .b(n1570), .O(n1576));
  andx g1276(.a(n1576), .b(pi120), .O(po045));
  andx g1277(.a(n1346), .b(n1553), .O(n1578));
  andx g1278(.a(n1349), .b(n1555), .O(n1579));
  andx g1279(.a(n1351), .b(pi105), .O(n1580));
  andx g1280(.a(n1353), .b(pi103), .O(n1581));
  orx  g1281(.a(n1581), .b(n1580), .O(n1582));
  orx  g1282(.a(n1582), .b(n1579), .O(n1583));
  orx  g1283(.a(n1583), .b(n1578), .O(po046));
  andx g1284(.a(n1179), .b(n458), .O(n1585));
  andx g1285(.a(n1201), .b(n500), .O(n1586));
  andx g1286(.a(n502), .b(pi134), .O(n1587));
  andx g1287(.a(n504), .b(pi135), .O(n1588));
  orx  g1288(.a(n1588), .b(n1587), .O(n1589));
  orx  g1289(.a(n1589), .b(n1586), .O(n1590));
  orx  g1290(.a(n1590), .b(n1585), .O(n1591));
  andx g1291(.a(n1591), .b(pi120), .O(po048));
  invx g1292(.a(n458), .O(n1593));
  orx  g1293(.a(n800), .b(n1593), .O(n1594));
  invx g1294(.a(n500), .O(n1595));
  orx  g1295(.a(n1081), .b(n1595), .O(n1596));
  invx g1296(.a(n502), .O(n1597));
  orx  g1297(.a(n1597), .b(n1086), .O(n1598));
  invx g1298(.a(n504), .O(n1599));
  orx  g1299(.a(n1599), .b(n1090), .O(n1600));
  andx g1300(.a(n1600), .b(n1598), .O(n1601));
  andx g1301(.a(n1601), .b(n1596), .O(n1602));
  andx g1302(.a(n1602), .b(n1594), .O(n1603));
  orx  g1303(.a(n1603), .b(n510), .O(po049));
  invx g1304(.a(pi174), .O(n1605));
  orx  g1305(.a(po071), .b(n1605), .O(po050));
  andx g1306(.a(n1464), .b(n802), .O(n1607));
  andx g1307(.a(n1474), .b(n1083), .O(n1608));
  andx g1308(.a(n1087), .b(pi142), .O(n1609));
  andx g1309(.a(n1091), .b(pi143), .O(n1610));
  orx  g1310(.a(n1610), .b(n1609), .O(n1611));
  orx  g1311(.a(n1611), .b(n1608), .O(n1612));
  orx  g1312(.a(n1612), .b(n1607), .O(n1613));
  andx g1313(.a(n1613), .b(pi120), .O(po054));
  invx g1314(.a(pi148), .O(n1615));
  andx g1315(.a(pi149), .b(n1615), .O(po055));
  invx g1316(.a(n1436), .O(po056));
  orx  g1317(.a(pi093), .b(pi064), .O(n1618));
  andx g1318(.a(n1618), .b(pi079), .O(n1619));
  orx  g1319(.a(n1619), .b(n795), .O(n1620));
  orx  g1320(.a(n1620), .b(n668), .O(po057));
  orx  g1321(.a(n1165), .b(n542), .O(n1622));
  andx g1322(.a(n1622), .b(n1167), .O(n1623));
  andx g1323(.a(n1623), .b(n420), .O(n1624));
  invx g1324(.a(n1624), .O(n1625));
  andx g1325(.a(n437), .b(pi089), .O(n1626));
  invx g1326(.a(n1626), .O(n1627));
  andx g1327(.a(pi007), .b(pi018), .O(n1628));
  andx g1328(.a(pi005), .b(n346), .O(n1629));
  orx  g1329(.a(n1629), .b(pi017), .O(n1630));
  orx  g1330(.a(n1630), .b(n1628), .O(n1631));
  andx g1331(.a(n446), .b(pi018), .O(n1632));
  andx g1332(.a(n448), .b(n346), .O(n1633));
  orx  g1333(.a(n1633), .b(n353), .O(n1634));
  orx  g1334(.a(n1634), .b(n1632), .O(n1635));
  andx g1335(.a(n1635), .b(n1631), .O(n1636));
  orx  g1336(.a(n1636), .b(n441), .O(n1637));
  andx g1337(.a(n1637), .b(n1627), .O(n1638));
  andx g1338(.a(n1638), .b(n1625), .O(po094));
  invx g1339(.a(po094), .O(n1640));
  andx g1340(.a(n1640), .b(n802), .O(n1641));
  andx g1341(.a(n1185), .b(n821), .O(n1642));
  orx  g1342(.a(n1642), .b(n1187), .O(n1643));
  orx  g1343(.a(n1643), .b(n421), .O(n1644));
  andx g1344(.a(n437), .b(pi086), .O(n1645));
  invx g1345(.a(n1645), .O(n1646));
  orx  g1346(.a(n1512), .b(n441), .O(n1647));
  andx g1347(.a(n1647), .b(n1646), .O(n1648));
  andx g1348(.a(n1648), .b(n1644), .O(po111));
  invx g1349(.a(po111), .O(n1650));
  andx g1350(.a(n1650), .b(n1083), .O(n1651));
  andx g1351(.a(n1087), .b(pi138), .O(n1652));
  andx g1352(.a(n1091), .b(pi139), .O(n1653));
  orx  g1353(.a(n1653), .b(n1652), .O(n1654));
  orx  g1354(.a(n1654), .b(n1651), .O(n1655));
  orx  g1355(.a(n1655), .b(n1641), .O(n1656));
  andx g1356(.a(n1656), .b(pi120), .O(po060));
  andx g1357(.a(n1118), .b(n458), .O(n1658));
  andx g1358(.a(n1145), .b(n500), .O(n1659));
  andx g1359(.a(n502), .b(pi132), .O(n1660));
  andx g1360(.a(n504), .b(pi133), .O(n1661));
  orx  g1361(.a(n1661), .b(n1660), .O(n1662));
  orx  g1362(.a(n1662), .b(n1659), .O(n1663));
  orx  g1363(.a(n1663), .b(n1658), .O(n1664));
  andx g1364(.a(n1664), .b(pi120), .O(po061));
  andx g1365(.a(n802), .b(n456), .O(n1666));
  andx g1366(.a(n1083), .b(n498), .O(n1667));
  andx g1367(.a(n1087), .b(pi129), .O(n1668));
  andx g1368(.a(n1091), .b(pi128), .O(n1669));
  orx  g1369(.a(n1669), .b(n1668), .O(n1670));
  orx  g1370(.a(n1670), .b(n1667), .O(n1671));
  orx  g1371(.a(n1671), .b(n1666), .O(n1672));
  andx g1372(.a(n1672), .b(pi120), .O(po062));
  andx g1373(.a(n1640), .b(n1346), .O(n1674));
  andx g1374(.a(n1650), .b(n1349), .O(n1675));
  andx g1375(.a(n1351), .b(pi100), .O(n1676));
  andx g1376(.a(n1353), .b(pi099), .O(n1677));
  orx  g1377(.a(n1677), .b(n1676), .O(n1678));
  orx  g1378(.a(n1678), .b(n1675), .O(n1679));
  orx  g1379(.a(n1679), .b(n1674), .O(po063));
  andx g1380(.a(pi058), .b(n925), .O(n1681));
  andx g1381(.a(n917), .b(pi065), .O(n1682));
  orx  g1382(.a(n1682), .b(n1681), .O(n1683));
  invx g1383(.a(n1683), .O(n1684));
  andx g1384(.a(pi042), .b(pi041), .O(n1685));
  andx g1385(.a(n828), .b(n463), .O(n1686));
  orx  g1386(.a(n1686), .b(n1685), .O(n1687));
  andx g1387(.a(n1687), .b(n812), .O(n1688));
  invx g1388(.a(n1688), .O(n1689));
  orx  g1389(.a(n1687), .b(n812), .O(n1690));
  andx g1390(.a(n1690), .b(n1689), .O(n1691));
  invx g1391(.a(n1691), .O(n1692));
  andx g1392(.a(n1692), .b(n1684), .O(n1693));
  andx g1393(.a(n1691), .b(n1683), .O(n1694));
  orx  g1394(.a(n1694), .b(n1693), .O(n1695));
  andx g1395(.a(pi067), .b(pi045), .O(n1696));
  invx g1396(.a(pi067), .O(n1697));
  andx g1397(.a(n1697), .b(n474), .O(n1698));
  orx  g1398(.a(n1698), .b(n1696), .O(n1699));
  invx g1399(.a(n1699), .O(n1700));
  andx g1400(.a(pi057), .b(pi059), .O(n1701));
  andx g1401(.a(n904), .b(n898), .O(n1702));
  orx  g1402(.a(n1702), .b(n1701), .O(n1703));
  andx g1403(.a(n1703), .b(n1700), .O(n1704));
  invx g1404(.a(n1704), .O(n1705));
  orx  g1405(.a(n1703), .b(n1700), .O(n1706));
  andx g1406(.a(n1706), .b(n1705), .O(n1707));
  invx g1407(.a(n1707), .O(n1708));
  andx g1408(.a(n1708), .b(n1695), .O(n1709));
  invx g1409(.a(n1709), .O(n1710));
  orx  g1410(.a(n1708), .b(n1695), .O(n1711));
  andx g1411(.a(n1711), .b(n1710), .O(po065));
  andx g1412(.a(pi036), .b(n383), .O(n1713));
  andx g1413(.a(n397), .b(pi015), .O(n1714));
  orx  g1414(.a(n1714), .b(n1713), .O(n1715));
  invx g1415(.a(n1715), .O(n1716));
  andx g1416(.a(pi027), .b(pi024), .O(n1717));
  andx g1417(.a(n312), .b(n671), .O(n1718));
  orx  g1418(.a(n1718), .b(n1717), .O(n1719));
  andx g1419(.a(n1719), .b(n346), .O(n1720));
  invx g1420(.a(n1720), .O(n1721));
  orx  g1421(.a(n1719), .b(n346), .O(n1722));
  andx g1422(.a(n1722), .b(n1721), .O(n1723));
  invx g1423(.a(n1723), .O(n1724));
  andx g1424(.a(n1724), .b(n1716), .O(n1725));
  andx g1425(.a(n1723), .b(n1715), .O(n1726));
  orx  g1426(.a(n1726), .b(n1725), .O(n1727));
  andx g1427(.a(pi006), .b(pi030), .O(n1728));
  invx g1428(.a(n1728), .O(n1729));
  orx  g1429(.a(pi006), .b(pi030), .O(n1730));
  andx g1430(.a(n1730), .b(n1729), .O(n1731));
  invx g1431(.a(n1731), .O(n1732));
  andx g1432(.a(n1732), .b(n335), .O(n1733));
  andx g1433(.a(n1731), .b(pi021), .O(n1734));
  orx  g1434(.a(n1734), .b(n1733), .O(n1735));
  invx g1435(.a(n1735), .O(n1736));
  andx g1436(.a(pi009), .b(pi012), .O(n1737));
  andx g1437(.a(n359), .b(n370), .O(n1738));
  orx  g1438(.a(n1738), .b(n1737), .O(n1739));
  andx g1439(.a(n1739), .b(n1736), .O(n1740));
  invx g1440(.a(n1740), .O(n1741));
  orx  g1441(.a(n1739), .b(n1736), .O(n1742));
  andx g1442(.a(n1742), .b(n1741), .O(n1743));
  invx g1443(.a(n1743), .O(n1744));
  andx g1444(.a(n1744), .b(n1727), .O(n1745));
  invx g1445(.a(n1745), .O(n1746));
  orx  g1446(.a(n1744), .b(n1727), .O(n1747));
  andx g1447(.a(n1747), .b(n1746), .O(n1748));
  invx g1448(.a(n1748), .O(po066));
  andx g1449(.a(n1424), .b(n458), .O(n1750));
  andx g1450(.a(n1436), .b(n500), .O(n1751));
  andx g1451(.a(n502), .b(pi116), .O(n1752));
  andx g1452(.a(n504), .b(pi115), .O(n1753));
  orx  g1453(.a(n1753), .b(n1752), .O(n1754));
  orx  g1454(.a(n1754), .b(n1751), .O(n1755));
  orx  g1455(.a(n1755), .b(n1750), .O(n1756));
  andx g1456(.a(n1756), .b(pi120), .O(po067));
  andx g1457(.a(n1346), .b(n1179), .O(n1758));
  andx g1458(.a(n1349), .b(n1201), .O(n1759));
  andx g1459(.a(n1351), .b(pi104), .O(n1760));
  andx g1460(.a(n1353), .b(pi108), .O(n1761));
  orx  g1461(.a(n1761), .b(n1760), .O(n1762));
  orx  g1462(.a(n1762), .b(n1759), .O(n1763));
  orx  g1463(.a(n1763), .b(n1758), .O(po068));
  andx g1464(.a(pi163), .b(pi159), .O(n1765));
  andx g1465(.a(pi162), .b(n1211), .O(n1766));
  orx  g1466(.a(n1766), .b(n1765), .O(n1767));
  orx  g1467(.a(n1767), .b(po071), .O(n1768));
  andx g1468(.a(n1768), .b(pi160), .O(po070));
  orx  g1469(.a(pi094), .b(pi064), .O(n1770));
  andx g1470(.a(n1770), .b(pi079), .O(n1771));
  orx  g1471(.a(n1771), .b(n1076), .O(n1772));
  orx  g1472(.a(n1772), .b(n977), .O(po072));
  invx g1473(.a(n1278), .O(po073));
  andx g1474(.a(n1346), .b(n1336), .O(n1775));
  andx g1475(.a(n1349), .b(n1338), .O(n1776));
  andx g1476(.a(n1351), .b(pi110), .O(n1777));
  andx g1477(.a(n1353), .b(pi102), .O(n1778));
  orx  g1478(.a(n1778), .b(n1777), .O(n1779));
  orx  g1479(.a(n1779), .b(n1776), .O(n1780));
  orx  g1480(.a(n1780), .b(n1775), .O(po075));
  invx g1481(.a(n1179), .O(po076));
  invx g1482(.a(n1196), .O(po077));
  andx g1483(.a(pi161), .b(pi160), .O(po078));
  andx g1484(.a(n1640), .b(n458), .O(n1785));
  andx g1485(.a(n1650), .b(n500), .O(n1786));
  andx g1486(.a(n502), .b(pi138), .O(n1787));
  andx g1487(.a(n504), .b(pi139), .O(n1788));
  orx  g1488(.a(n1788), .b(n1787), .O(n1789));
  orx  g1489(.a(n1789), .b(n1786), .O(n1790));
  orx  g1490(.a(n1790), .b(n1785), .O(n1791));
  andx g1491(.a(n1791), .b(pi120), .O(po079));
  andx g1492(.a(n1346), .b(n1278), .O(n1793));
  andx g1493(.a(n1349), .b(n1290), .O(n1794));
  andx g1494(.a(n1351), .b(pi111), .O(n1795));
  andx g1495(.a(n1353), .b(pi112), .O(n1796));
  orx  g1496(.a(n1796), .b(n1795), .O(n1797));
  orx  g1497(.a(n1797), .b(n1794), .O(n1798));
  orx  g1498(.a(n1798), .b(n1793), .O(po080));
  andx g1499(.a(n1527), .b(n458), .O(n1800));
  andx g1500(.a(n1540), .b(n500), .O(n1801));
  andx g1501(.a(n502), .b(pi140), .O(n1802));
  andx g1502(.a(n504), .b(pi141), .O(n1803));
  orx  g1503(.a(n1803), .b(n1802), .O(n1804));
  orx  g1504(.a(n1804), .b(n1801), .O(n1805));
  orx  g1505(.a(n1805), .b(n1800), .O(n1806));
  andx g1506(.a(n1806), .b(pi120), .O(po084));
  andx g1507(.a(n1527), .b(n802), .O(n1808));
  andx g1508(.a(n1540), .b(n1083), .O(n1809));
  andx g1509(.a(n1087), .b(pi140), .O(n1810));
  andx g1510(.a(n1091), .b(pi141), .O(n1811));
  orx  g1511(.a(n1811), .b(n1810), .O(n1812));
  orx  g1512(.a(n1812), .b(n1809), .O(n1813));
  orx  g1513(.a(n1813), .b(n1808), .O(n1814));
  andx g1514(.a(n1814), .b(pi120), .O(po085));
  andx g1515(.a(pi164), .b(pi159), .O(n1816));
  andx g1516(.a(pi165), .b(n1211), .O(n1817));
  orx  g1517(.a(n1817), .b(n1816), .O(n1818));
  orx  g1518(.a(n1818), .b(po071), .O(n1819));
  andx g1519(.a(n1819), .b(pi160), .O(po086));
  andx g1520(.a(n1306), .b(n1278), .O(n1821));
  andx g1521(.a(n1309), .b(n1290), .O(n1822));
  andx g1522(.a(n1311), .b(pi111), .O(n1823));
  andx g1523(.a(n1313), .b(pi112), .O(n1824));
  orx  g1524(.a(n1824), .b(n1823), .O(n1825));
  orx  g1525(.a(n1825), .b(n1822), .O(n1826));
  orx  g1526(.a(n1826), .b(n1821), .O(po087));
  andx g1527(.a(n1346), .b(n1527), .O(n1828));
  andx g1528(.a(n1540), .b(n1349), .O(n1829));
  andx g1529(.a(n1351), .b(pi107), .O(n1830));
  andx g1530(.a(n1353), .b(pi106), .O(n1831));
  orx  g1531(.a(n1831), .b(n1830), .O(n1832));
  orx  g1532(.a(n1832), .b(n1829), .O(n1833));
  orx  g1533(.a(n1833), .b(n1828), .O(po088));
  invx g1534(.a(pi171), .O(po089));
  andx g1535(.a(n1640), .b(n1306), .O(n1836));
  andx g1536(.a(n1650), .b(n1309), .O(n1837));
  andx g1537(.a(n1311), .b(pi100), .O(n1838));
  andx g1538(.a(n1313), .b(pi099), .O(n1839));
  orx  g1539(.a(n1839), .b(n1838), .O(n1840));
  orx  g1540(.a(n1840), .b(n1837), .O(n1841));
  orx  g1541(.a(n1841), .b(n1836), .O(po091));
  invx g1542(.a(n1474), .O(po092));
  orx  g1543(.a(pi156), .b(n1214), .O(po093));
  invx g1544(.a(n1469), .O(n1845));
  andx g1545(.a(n1181), .b(n866), .O(n1846));
  andx g1546(.a(n1846), .b(n1643), .O(n1847));
  andx g1547(.a(n1847), .b(n1283), .O(n1848));
  andx g1548(.a(n1848), .b(n1533), .O(n1849));
  andx g1549(.a(n1849), .b(po077), .O(n1850));
  andx g1550(.a(n1850), .b(n1845), .O(po095));
  invx g1551(.a(n1464), .O(po096));
  andx g1552(.a(pi166), .b(pi159), .O(n1853));
  andx g1553(.a(pi167), .b(n1211), .O(n1854));
  orx  g1554(.a(n1854), .b(n1853), .O(n1855));
  orx  g1555(.a(n1855), .b(po071), .O(n1856));
  andx g1556(.a(n1856), .b(pi160), .O(po097));
  andx g1557(.a(n1464), .b(n1306), .O(n1858));
  andx g1558(.a(n1474), .b(n1309), .O(n1859));
  andx g1559(.a(n1311), .b(pi098), .O(n1860));
  andx g1560(.a(n1313), .b(pi109), .O(n1861));
  orx  g1561(.a(n1861), .b(n1860), .O(n1862));
  orx  g1562(.a(n1862), .b(n1859), .O(n1863));
  orx  g1563(.a(n1863), .b(n1858), .O(po101));
  andx g1564(.a(n849), .b(n810), .O(n1865));
  andx g1565(.a(n852), .b(n817), .O(n1866));
  orx  g1566(.a(n1866), .b(n1865), .O(n1867));
  invx g1567(.a(n1867), .O(n1868));
  andx g1568(.a(n1697), .b(n464), .O(n1869));
  invx g1569(.a(n1869), .O(n1870));
  orx  g1570(.a(pi068), .b(n464), .O(n1871));
  andx g1571(.a(n1871), .b(n1870), .O(n1872));
  andx g1572(.a(n1872), .b(n476), .O(n1873));
  invx g1573(.a(n1873), .O(n1874));
  orx  g1574(.a(n1872), .b(n476), .O(n1875));
  andx g1575(.a(n1875), .b(n1874), .O(n1876));
  andx g1576(.a(n1876), .b(n466), .O(n1877));
  invx g1577(.a(n1877), .O(n1878));
  orx  g1578(.a(n1876), .b(n466), .O(n1879));
  andx g1579(.a(n1879), .b(n1878), .O(n1880));
  invx g1580(.a(n1880), .O(n1881));
  andx g1581(.a(n1881), .b(n830), .O(n1882));
  andx g1582(.a(n1880), .b(n831), .O(n1883));
  orx  g1583(.a(n1883), .b(n1882), .O(n1884));
  andx g1584(.a(n1884), .b(n1868), .O(n1885));
  invx g1585(.a(n1885), .O(n1886));
  orx  g1586(.a(n1884), .b(n1868), .O(n1887));
  andx g1587(.a(n1887), .b(n1886), .O(n1888));
  invx g1588(.a(n1888), .O(n1889));
  andx g1589(.a(n907), .b(n910), .O(n1890));
  andx g1590(.a(n938), .b(n901), .O(n1891));
  orx  g1591(.a(n1891), .b(n1890), .O(n1892));
  invx g1592(.a(n1892), .O(n1893));
  andx g1593(.a(n1893), .b(n932), .O(n1894));
  andx g1594(.a(n1892), .b(n933), .O(n1895));
  orx  g1595(.a(n1895), .b(n1894), .O(n1896));
  andx g1596(.a(n1896), .b(n1889), .O(n1897));
  invx g1597(.a(n1897), .O(n1898));
  orx  g1598(.a(n1896), .b(n1889), .O(n1899));
  andx g1599(.a(n1899), .b(n1898), .O(po122));
  invx g1600(.a(po122), .O(n1901));
  invx g1601(.a(po065), .O(n1902));
  andx g1602(.a(pi171), .b(pi170), .O(po115));
  andx g1603(.a(pi173), .b(pi172), .O(n1904));
  andx g1604(.a(pi151), .b(pi150), .O(n1905));
  andx g1605(.a(n1905), .b(n1904), .O(n1906));
  andx g1606(.a(n1906), .b(po115), .O(n1907));
  andx g1607(.a(n1907), .b(n1748), .O(n1908));
  andx g1608(.a(n1908), .b(n1902), .O(n1909));
  andx g1609(.a(n1909), .b(n1396), .O(n1910));
  andx g1610(.a(n1910), .b(n1901), .O(po102));
  andx g1611(.a(n1424), .b(n1306), .O(n1912));
  andx g1612(.a(n1436), .b(n1309), .O(n1913));
  andx g1613(.a(n1311), .b(pi113), .O(n1914));
  andx g1614(.a(n1313), .b(pi114), .O(n1915));
  orx  g1615(.a(n1915), .b(n1914), .O(n1916));
  orx  g1616(.a(n1916), .b(n1913), .O(n1917));
  orx  g1617(.a(n1917), .b(n1912), .O(po106));
  andx g1618(.a(n1460), .b(n1254), .O(n1919));
  andx g1619(.a(n1919), .b(n748), .O(n1920));
  andx g1620(.a(n1636), .b(n452), .O(n1921));
  andx g1621(.a(n1420), .b(n1332), .O(n1922));
  andx g1622(.a(n1274), .b(n1114), .O(n1923));
  andx g1623(.a(n1923), .b(n1922), .O(n1924));
  andx g1624(.a(n1924), .b(n1921), .O(n1925));
  andx g1625(.a(n1925), .b(n1920), .O(po107));
  invx g1626(.a(n1201), .O(po108));
  invx g1627(.a(pi151), .O(po109));
  andx g1628(.a(n1468), .b(pi069), .O(n1929));
  andx g1629(.a(n1467), .b(n1226), .O(n1930));
  orx  g1630(.a(n1930), .b(n1929), .O(po110));
  invx g1631(.a(pi150), .O(po112));
  invx g1632(.a(n1448), .O(n1933));
  invx g1633(.a(n1623), .O(n1934));
  invx g1634(.a(n1319), .O(n1935));
  andx g1635(.a(n1935), .b(n434), .O(n1936));
  andx g1636(.a(n1936), .b(n1102), .O(n1937));
  andx g1637(.a(n1937), .b(n1408), .O(n1938));
  andx g1638(.a(n1938), .b(n1934), .O(n1939));
  andx g1639(.a(n1939), .b(n1242), .O(n1940));
  andx g1640(.a(n1940), .b(n1933), .O(n1941));
  invx g1641(.a(n1174), .O(n1942));
  invx g1642(.a(n1262), .O(n1943));
  andx g1643(.a(n1943), .b(n1942), .O(n1944));
  andx g1644(.a(n1944), .b(n1941), .O(po114));
  andx g1645(.a(pi168), .b(pi159), .O(n1946));
  andx g1646(.a(pi169), .b(n1211), .O(n1947));
  orx  g1647(.a(n1947), .b(n1946), .O(n1948));
  orx  g1648(.a(n1948), .b(po071), .O(n1949));
  andx g1649(.a(n1949), .b(pi160), .O(po116));
  andx g1650(.a(n1464), .b(n458), .O(n1951));
  andx g1651(.a(n1474), .b(n500), .O(n1952));
  andx g1652(.a(n502), .b(pi142), .O(n1953));
  andx g1653(.a(n504), .b(pi143), .O(n1954));
  orx  g1654(.a(n1954), .b(n1953), .O(n1955));
  orx  g1655(.a(n1955), .b(n1952), .O(n1956));
  orx  g1656(.a(n1956), .b(n1951), .O(n1957));
  andx g1657(.a(n1957), .b(pi120), .O(po117));
  invx g1658(.a(pi175), .O(n1959));
  orx  g1659(.a(po071), .b(n1959), .O(po118));
  andx g1660(.a(n1306), .b(n456), .O(n1961));
  andx g1661(.a(n1309), .b(n498), .O(n1962));
  andx g1662(.a(n1311), .b(pi096), .O(n1963));
  andx g1663(.a(n1313), .b(pi097), .O(n1964));
  orx  g1664(.a(n1964), .b(n1963), .O(n1965));
  orx  g1665(.a(n1965), .b(n1962), .O(n1966));
  orx  g1666(.a(n1966), .b(n1961), .O(po119));
  invx g1667(.a(n1904), .O(po121));
  bufx g1668(.a(pi148), .O(po012));
  invx g1669(.a(pi177), .O(po026));
  bufx g1670(.a(pi146), .O(po027));
  orx  g1671(.a(n1158), .b(n1155), .O(po028));
  bufx g1672(.a(pi176), .O(po029));
  bufx g1673(.a(pi146), .O(po030));
  bufx g1674(.a(pi146), .O(po037));
  invx g1675(.a(pi177), .O(po047));
  bufx g1676(.a(pi146), .O(po053));
  bufx g1677(.a(pi120), .O(po058));
  orx  g1678(.a(n416), .b(n407), .O(po059));
  bufx g1679(.a(pi065), .O(po069));
  invx g1680(.a(pi176), .O(po074));
  andx g1681(.a(n1157), .b(n893), .O(po082));
  andx g1682(.a(n543), .b(n406), .O(po083));
  orx  g1683(.a(n1217), .b(n1210), .O(po090));
  bufx g1684(.a(pi066), .O(po098));
  bufx g1685(.a(pi160), .O(po099));
  bufx g1686(.a(pi160), .O(po100));
  bufx g1687(.a(pi066), .O(po104));
  bufx g1688(.a(pi146), .O(po113));
endmodule


