// Benchmark "h264lut_coeff" written by ABC on Fri Feb  7 13:43:12 2014

module h264lut_coeff ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10;
  wire n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
    n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
    n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63,
    n64, n65, n66, n67, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n213, n214, n215, n217, n218,
    n219, n220, n221, n222, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710;
  bufx g000(.A(n632), .O(n21));
  invx g001(.A(n645), .O(n22));
  bufx g002(.A(n599), .O(n23));
  bufx g003(.A(n569), .O(n24));
  bufx g004(.A(n398), .O(n25));
  bufx g005(.A(n613), .O(n26));
  bufx g006(.A(n350), .O(n27));
  bufx g007(.A(n617), .O(n28));
  bufx g008(.A(n600), .O(n29));
  bufx g009(.A(n587), .O(n30));
  bufx g010(.A(n625), .O(n31));
  bufx g011(.A(n625), .O(n32));
  bufx g012(.A(n561), .O(n33));
  bufx g013(.A(n621), .O(n34));
  bufx g014(.A(n680), .O(n35));
  bufx g015(.A(n680), .O(n36));
  bufx g016(.A(n675), .O(n37));
  bufx g017(.A(n626), .O(n38));
  bufx g018(.A(n704), .O(n39));
  bufx g019(.A(n704), .O(n40));
  invx g020(.A(n650), .O(n41));
  invx g021(.A(n41), .O(n42));
  invx g022(.A(n41), .O(n43));
  bufx g023(.A(n667), .O(n44));
  bufx g024(.A(n709), .O(n45));
  bufx g025(.A(n669), .O(n46));
  bufx g026(.A(n391), .O(n47));
  bufx g027(.A(n620), .O(n48));
  bufx g028(.A(n657), .O(n49));
  bufx g029(.A(n657), .O(n50));
  bufx g030(.A(n651), .O(n51));
  bufx g031(.A(n651), .O(n52));
  bufx g032(.A(n603), .O(n53));
  bufx g033(.A(n674), .O(n54));
  bufx g034(.A(n624), .O(n55));
  bufx g035(.A(n604), .O(n56));
  bufx g036(.A(n506), .O(n57));
  bufx g037(.A(n646), .O(n58));
  bufx g038(.A(n646), .O(n59));
  bufx g039(.A(n415), .O(n60));
  bufx g040(.A(n415), .O(n61));
  orx  g041(.A(n66), .B(n63), .O(po10));
  andx g042(.A(n627), .B(n64), .O(n63));
  orx  g043(.A(n65), .B(n288), .O(n64));
  andx g044(.A(n652), .B(n589), .O(n65));
  andx g045(.A(n67), .B(pi0), .O(n66));
  andx g046(.A(n31), .B(n653), .O(n67));
  orx  g047(.A(n70), .B(n69), .O(po09));
  orx  g048(.A(n567), .B(n236), .O(n69));
  orx  g049(.A(n92), .B(n71), .O(n70));
  orx  g050(.A(n331), .B(n72), .O(n71));
  andx g051(.A(n43), .B(n73), .O(n72));
  orx  g052(.A(n506), .B(n29), .O(n73));
  andx g053(.A(n83), .B(n75), .O(po08));
  andx g054(.A(n79), .B(n76), .O(n75));
  invx g055(.A(n77), .O(n76));
  orx  g056(.A(n78), .B(n440), .O(n77));
  orx  g057(.A(n533), .B(n497), .O(n78));
  andx g058(.A(n81), .B(n80), .O(n79));
  orx  g059(.A(n369), .B(n655), .O(n80));
  andx g060(.A(n82), .B(n262), .O(n81));
  orx  g061(.A(n112), .B(n633), .O(n82));
  andx g062(.A(n89), .B(n84), .O(n83));
  andx g063(.A(n85), .B(n189), .O(n84));
  andx g064(.A(n87), .B(n86), .O(n85));
  orx  g065(.A(n605), .B(n368), .O(n86));
  invx g066(.A(n88), .O(n87));
  andx g067(.A(n48), .B(n24), .O(n88));
  invx g068(.A(n90), .O(n89));
  orx  g069(.A(n91), .B(n208), .O(n90));
  orx  g070(.A(n556), .B(n92), .O(n91));
  orx  g071(.A(n96), .B(n93), .O(n92));
  orx  g072(.A(n95), .B(n94), .O(n93));
  orx  g073(.A(n333), .B(n204), .O(n94));
  orx  g074(.A(n316), .B(n152), .O(n95));
  orx  g075(.A(n100), .B(n97), .O(n96));
  orx  g076(.A(n99), .B(n98), .O(n97));
  andx g077(.A(n38), .B(n35), .O(n98));
  andx g078(.A(n22), .B(n387), .O(n99));
  orx  g079(.A(n102), .B(n101), .O(n100));
  orx  g080(.A(n419), .B(n330), .O(n101));
  andx g081(.A(n665), .B(n29), .O(n102));
  andx g082(.A(n130), .B(n104), .O(po07));
  andx g083(.A(n117), .B(n105), .O(n104));
  andx g084(.A(n109), .B(n106), .O(n105));
  invx g085(.A(n107), .O(n106));
  orx  g086(.A(n108), .B(n427), .O(n107));
  orx  g087(.A(n483), .B(n533), .O(n108));
  andx g088(.A(n110), .B(n366), .O(n109));
  andx g089(.A(n113), .B(n111), .O(n110));
  orx  g090(.A(n605), .B(n112), .O(n111));
  invx g091(.A(n53), .O(n112));
  orx  g092(.A(n114), .B(n180), .O(n113));
  invx g093(.A(n115), .O(n114));
  orx  g094(.A(n116), .B(n54), .O(n115));
  orx  g095(.A(n649), .B(n595), .O(n116));
  andx g096(.A(n125), .B(n118), .O(n117));
  andx g097(.A(n122), .B(n119), .O(n118));
  orx  g098(.A(n121), .B(n120), .O(n119));
  invx g099(.A(n506), .O(n120));
  andx g100(.A(n379), .B(n44), .O(n121));
  andx g101(.A(n124), .B(n123), .O(n122));
  orx  g102(.A(n263), .B(n44), .O(n123));
  orx  g103(.A(n197), .B(n655), .O(n124));
  andx g104(.A(n129), .B(n126), .O(n125));
  orx  g105(.A(n127), .B(n380), .O(n126));
  andx g106(.A(n128), .B(n645), .O(n127));
  invx g107(.A(n54), .O(n128));
  orx  g108(.A(n193), .B(n505), .O(n129));
  andx g109(.A(n144), .B(n131), .O(n130));
  andx g110(.A(n137), .B(n132), .O(n131));
  invx g111(.A(n133), .O(n132));
  orx  g112(.A(n135), .B(n134), .O(n133));
  andx g113(.A(n457), .B(n604), .O(n134));
  orx  g114(.A(n136), .B(n558), .O(n135));
  andx g115(.A(n355), .B(n36), .O(n136));
  andx g116(.A(n140), .B(n138), .O(n137));
  invx g117(.A(n139), .O(n138));
  andx g118(.A(n32), .B(n654), .O(n139));
  andx g119(.A(n143), .B(n141), .O(n140));
  invx g120(.A(n142), .O(n141));
  andx g121(.A(n665), .B(n587), .O(n142));
  orx  g122(.A(n190), .B(n676), .O(n143));
  andx g123(.A(n150), .B(n145), .O(n144));
  andx g124(.A(n147), .B(n146), .O(n145));
  invx g125(.A(n336), .O(n146));
  andx g126(.A(n149), .B(n148), .O(n147));
  orx  g127(.A(n193), .B(n678), .O(n148));
  invx g128(.A(n239), .O(n149));
  invx g129(.A(n151), .O(n150));
  orx  g130(.A(n208), .B(n152), .O(n151));
  orx  g131(.A(n155), .B(n153), .O(n152));
  orx  g132(.A(n154), .B(n264), .O(n153));
  andx g133(.A(n26), .B(n47), .O(n154));
  orx  g134(.A(n442), .B(n156), .O(n155));
  orx  g135(.A(n498), .B(n526), .O(n156));
  andx g136(.A(n186), .B(n158), .O(po06));
  andx g137(.A(n171), .B(n159), .O(n158));
  andx g138(.A(n165), .B(n160), .O(n159));
  invx g139(.A(n161), .O(n160));
  orx  g140(.A(n164), .B(n162), .O(n161));
  andx g141(.A(n48), .B(n163), .O(n162));
  orx  g142(.A(n621), .B(n40), .O(n163));
  orx  g143(.A(n246), .B(n629), .O(n164));
  andx g144(.A(n168), .B(n166), .O(n165));
  orx  g145(.A(n167), .B(n678), .O(n166));
  andx g146(.A(n369), .B(n190), .O(n167));
  invx g147(.A(n169), .O(n168));
  andx g148(.A(n170), .B(n675), .O(n169));
  orx  g149(.A(n420), .B(n32), .O(n170));
  andx g150(.A(n182), .B(n172), .O(n171));
  andx g151(.A(n178), .B(n173), .O(n172));
  orx  g152(.A(n174), .B(n618), .O(n173));
  andx g153(.A(n176), .B(n175), .O(n174));
  andx g154(.A(n197), .B(n199), .O(n175));
  andx g155(.A(n177), .B(n263), .O(n176));
  invx g156(.A(n467), .O(n177));
  andx g157(.A(n181), .B(n179), .O(n178));
  orx  g158(.A(n384), .B(n180), .O(n179));
  invx g159(.A(n569), .O(n180));
  orx  g160(.A(n371), .B(n698), .O(n181));
  invx g161(.A(n183), .O(n182));
  orx  g162(.A(n185), .B(n184), .O(n183));
  andx g163(.A(n686), .B(n355), .O(n184));
  andx g164(.A(n25), .B(n680), .O(n185));
  andx g165(.A(n200), .B(n187), .O(n186));
  andx g166(.A(n195), .B(n188), .O(n187));
  andx g167(.A(n191), .B(n189), .O(n188));
  orx  g168(.A(n190), .B(n633), .O(n189));
  invx g169(.A(n626), .O(n190));
  andx g170(.A(n194), .B(n192), .O(n191));
  orx  g171(.A(n193), .B(n44), .O(n192));
  invx g172(.A(n47), .O(n193));
  invx g173(.A(n253), .O(n194));
  andx g174(.A(n198), .B(n196), .O(n195));
  orx  g175(.A(n197), .B(n605), .O(n196));
  invx g176(.A(n58), .O(n197));
  orx  g177(.A(n655), .B(n199), .O(n198));
  invx g178(.A(n33), .O(n199));
  invx g179(.A(n201), .O(n200));
  orx  g180(.A(n211), .B(n202), .O(n201));
  orx  g181(.A(n203), .B(n538), .O(n202));
  orx  g182(.A(n208), .B(n204), .O(n203));
  orx  g183(.A(n207), .B(n205), .O(n204));
  orx  g184(.A(n481), .B(n206), .O(n205));
  andx g185(.A(n51), .B(n598), .O(n206));
  andx g186(.A(n639), .B(n295), .O(n207));
  orx  g187(.A(n210), .B(n209), .O(n208));
  andx g188(.A(n42), .B(n27), .O(n209));
  andx g189(.A(n279), .B(n288), .O(n210));
  orx  g190(.A(n310), .B(n430), .O(n211));
  orx  g191(.A(n214), .B(n213), .O(po05));
  orx  g192(.A(n218), .B(n231), .O(n213));
  orx  g193(.A(n413), .B(n215), .O(n214));
  andx g194(.A(n22), .B(n60), .O(n215));
  orx  g195(.A(n221), .B(n217), .O(po04));
  orx  g196(.A(n218), .B(n229), .O(n217));
  orx  g197(.A(n268), .B(n219), .O(n218));
  orx  g198(.A(n410), .B(n220), .O(n219));
  andx g199(.A(n26), .B(n61), .O(n220));
  orx  g200(.A(n406), .B(n222), .O(n221));
  andx g201(.A(n677), .B(n60), .O(n222));
  orx  g202(.A(n275), .B(n224), .O(po03));
  orx  g203(.A(n233), .B(n225), .O(n224));
  orx  g204(.A(n227), .B(n226), .O(n225));
  orx  g205(.A(n306), .B(n425), .O(n226));
  orx  g206(.A(n536), .B(n228), .O(n227));
  orx  g207(.A(n231), .B(n229), .O(n228));
  orx  g208(.A(n230), .B(n407), .O(n229));
  andx g209(.A(n666), .B(n61), .O(n230));
  orx  g210(.A(n232), .B(n409), .O(n231));
  andx g211(.A(n687), .B(n60), .O(n232));
  orx  g212(.A(n270), .B(n234), .O(n233));
  orx  g213(.A(n268), .B(n235), .O(n234));
  orx  g214(.A(n264), .B(n236), .O(n235));
  orx  g215(.A(n254), .B(n237), .O(n236));
  orx  g216(.A(n251), .B(n238), .O(n237));
  orx  g217(.A(n250), .B(n239), .O(n238));
  orx  g218(.A(n247), .B(n240), .O(n239));
  orx  g219(.A(n244), .B(n241), .O(n240));
  orx  g220(.A(n243), .B(n242), .O(n241));
  andx g221(.A(n36), .B(n31), .O(n242));
  andx g222(.A(n521), .B(n383), .O(n243));
  orx  g223(.A(n246), .B(n245), .O(n244));
  andx g224(.A(n46), .B(n27), .O(n245));
  andx g225(.A(n29), .B(n48), .O(n246));
  orx  g226(.A(n249), .B(n248), .O(n247));
  orx  g227(.A(n484), .B(n440), .O(n248));
  orx  g228(.A(n497), .B(n495), .O(n249));
  andx g229(.A(n57), .B(n26), .O(n250));
  orx  g230(.A(n253), .B(n252), .O(n251));
  andx g231(.A(n685), .B(n279), .O(n252));
  andx g232(.A(n29), .B(n52), .O(n253));
  orx  g233(.A(n259), .B(n255), .O(n254));
  orx  g234(.A(n257), .B(n256), .O(n255));
  andx g235(.A(n34), .B(n612), .O(n256));
  andx g236(.A(n24), .B(n258), .O(n257));
  orx  g237(.A(n42), .B(n48), .O(n258));
  orx  g238(.A(n261), .B(n260), .O(n259));
  orx  g239(.A(n566), .B(n446), .O(n260));
  invx g240(.A(n262), .O(n261));
  orx  g241(.A(n263), .B(n645), .O(n262));
  invx g242(.A(n601), .O(n263));
  orx  g243(.A(n266), .B(n265), .O(n264));
  andx g244(.A(n686), .B(n295), .O(n265));
  andx g245(.A(n697), .B(n267), .O(n266));
  orx  g246(.A(n40), .B(n598), .O(n267));
  orx  g247(.A(n269), .B(n414), .O(n268));
  andx g248(.A(n52), .B(n61), .O(n269));
  orx  g249(.A(n274), .B(n271), .O(n270));
  orx  g250(.A(n273), .B(n272), .O(n271));
  andx g251(.A(n666), .B(n49), .O(n272));
  andx g252(.A(n35), .B(n24), .O(n273));
  andx g253(.A(n40), .B(n644), .O(n274));
  orx  g254(.A(n289), .B(n276), .O(n275));
  orx  g255(.A(n281), .B(n277), .O(n276));
  orx  g256(.A(n280), .B(n278), .O(n277));
  andx g257(.A(n42), .B(n279), .O(n278));
  orx  g258(.A(n506), .B(n27), .O(n279));
  andx g259(.A(n46), .B(n29), .O(n280));
  orx  g260(.A(n287), .B(n282), .O(n281));
  orx  g261(.A(n284), .B(n283), .O(n282));
  andx g262(.A(n586), .B(n47), .O(n283));
  andx g263(.A(n28), .B(n285), .O(n284));
  orx  g264(.A(n60), .B(n286), .O(n285));
  orx  g265(.A(n58), .B(n601), .O(n286));
  andx g266(.A(n57), .B(n288), .O(n287));
  orx  g267(.A(n640), .B(n52), .O(n288));
  orx  g268(.A(n299), .B(n290), .O(n289));
  orx  g269(.A(n297), .B(n291), .O(n290));
  orx  g270(.A(n294), .B(n292), .O(n291));
  andx g271(.A(n30), .B(n293), .O(n292));
  orx  g272(.A(n697), .B(n612), .O(n293));
  andx g273(.A(n296), .B(n295), .O(n294));
  orx  g274(.A(n59), .B(n47), .O(n295));
  orx  g275(.A(n677), .B(n363), .O(n296));
  andx g276(.A(n51), .B(n298), .O(n297));
  orx  g277(.A(n38), .B(n23), .O(n298));
  orx  g278(.A(n402), .B(n300), .O(n299));
  orx  g279(.A(n533), .B(n324), .O(n300));
  orx  g280(.A(n373), .B(n302), .O(po02));
  orx  g281(.A(n346), .B(n303), .O(n302));
  orx  g282(.A(n339), .B(n304), .O(n303));
  orx  g283(.A(n309), .B(n305), .O(n304));
  orx  g284(.A(n306), .B(n529), .O(n305));
  orx  g285(.A(n308), .B(n307), .O(n306));
  andx g286(.A(n37), .B(n59), .O(n307));
  andx g287(.A(n28), .B(n47), .O(n308));
  orx  g288(.A(n333), .B(n310), .O(n309));
  orx  g289(.A(n321), .B(n311), .O(n310));
  orx  g290(.A(n314), .B(n312), .O(n311));
  orx  g291(.A(n548), .B(n313), .O(n312));
  orx  g292(.A(n445), .B(n492), .O(n313));
  orx  g293(.A(n318), .B(n315), .O(n314));
  orx  g294(.A(n317), .B(n316), .O(n315));
  andx g295(.A(n46), .B(n57), .O(n316));
  andx g296(.A(n21), .B(n32), .O(n317));
  orx  g297(.A(n320), .B(n319), .O(n318));
  andx g298(.A(n30), .B(n644), .O(n319));
  andx g299(.A(n37), .B(n25), .O(n320));
  orx  g300(.A(n328), .B(n322), .O(n321));
  orx  g301(.A(n325), .B(n323), .O(n322));
  orx  g302(.A(n324), .B(n427), .O(n323));
  andx g303(.A(n457), .B(n35), .O(n324));
  andx g304(.A(n56), .B(n326), .O(n325));
  orx  g305(.A(n626), .B(n327), .O(n326));
  orx  g306(.A(n33), .B(n39), .O(n327));
  orx  g307(.A(n332), .B(n329), .O(n328));
  orx  g308(.A(n331), .B(n330), .O(n329));
  andx g309(.A(n420), .B(n36), .O(n330));
  andx g310(.A(n383), .B(n640), .O(n331));
  orx  g311(.A(n526), .B(n566), .O(n332));
  orx  g312(.A(n336), .B(n334), .O(n333));
  orx  g313(.A(n483), .B(n335), .O(n334));
  andx g314(.A(n54), .B(n27), .O(n335));
  orx  g315(.A(n338), .B(n337), .O(n336));
  andx g316(.A(n677), .B(n50), .O(n337));
  andx g317(.A(n35), .B(n600), .O(n338));
  orx  g318(.A(n343), .B(n340), .O(n339));
  orx  g319(.A(n342), .B(n341), .O(n340));
  andx g320(.A(n39), .B(n691), .O(n341));
  andx g321(.A(n52), .B(n59), .O(n342));
  orx  g322(.A(n345), .B(n344), .O(n343));
  andx g323(.A(n617), .B(n49), .O(n344));
  andx g324(.A(n30), .B(n26), .O(n345));
  orx  g325(.A(n356), .B(n347), .O(n346));
  orx  g326(.A(n352), .B(n348), .O(n347));
  orx  g327(.A(n351), .B(n349), .O(n348));
  andx g328(.A(n640), .B(n27), .O(n349));
  orx  g329(.A(n621), .B(n55), .O(n350));
  andx g330(.A(n36), .B(n624), .O(n351));
  orx  g331(.A(n354), .B(n353), .O(n352));
  andx g332(.A(n677), .B(n25), .O(n353));
  andx g333(.A(n355), .B(n48), .O(n354));
  orx  g334(.A(n587), .B(n57), .O(n355));
  orx  g335(.A(n364), .B(n357), .O(n356));
  orx  g336(.A(n362), .B(n358), .O(n357));
  andx g337(.A(n56), .B(n359), .O(n358));
  orx  g338(.A(n361), .B(n360), .O(n359));
  orx  g339(.A(n53), .B(n416), .O(n360));
  orx  g340(.A(n599), .B(n50), .O(n361));
  andx g341(.A(n38), .B(n363), .O(n362));
  orx  g342(.A(n650), .B(n666), .O(n363));
  invx g343(.A(n365), .O(n364));
  andx g344(.A(n370), .B(n366), .O(n365));
  orx  g345(.A(n41), .B(n367), .O(n366));
  andx g346(.A(n369), .B(n368), .O(n367));
  invx g347(.A(n602), .O(n368));
  invx g348(.A(n49), .O(n369));
  orx  g349(.A(n688), .B(n371), .O(n370));
  invx g350(.A(n372), .O(n371));
  orx  g351(.A(n599), .B(n55), .O(n372));
  orx  g352(.A(n403), .B(n374), .O(n373));
  orx  g353(.A(n392), .B(n375), .O(n374));
  orx  g354(.A(n385), .B(n376), .O(n375));
  invx g355(.A(n377), .O(n376));
  andx g356(.A(n381), .B(n378), .O(n377));
  orx  g357(.A(n380), .B(n379), .O(n378));
  andx g358(.A(n698), .B(n618), .O(n379));
  invx g359(.A(n621), .O(n380));
  orx  g360(.A(n384), .B(n382), .O(n381));
  invx g361(.A(n383), .O(n382));
  orx  g362(.A(n569), .B(n29), .O(n383));
  andx g363(.A(n692), .B(n44), .O(n384));
  orx  g364(.A(n388), .B(n386), .O(n385));
  andx g365(.A(n387), .B(n612), .O(n386));
  orx  g366(.A(n569), .B(n57), .O(n387));
  andx g367(.A(n669), .B(n389), .O(n388));
  orx  g368(.A(n25), .B(n390), .O(n389));
  orx  g369(.A(n621), .B(n47), .O(n390));
  orx  g370(.A(n587), .B(n457), .O(n391));
  orx  g371(.A(n399), .B(n393), .O(n392));
  orx  g372(.A(n396), .B(n394), .O(n393));
  andx g373(.A(n57), .B(n395), .O(n394));
  orx  g374(.A(n52), .B(n677), .O(n395));
  andx g375(.A(n697), .B(n397), .O(n396));
  orx  g376(.A(n591), .B(n25), .O(n397));
  orx  g377(.A(n569), .B(n601), .O(n398));
  orx  g378(.A(n402), .B(n400), .O(n399));
  andx g379(.A(n23), .B(n401), .O(n400));
  orx  g380(.A(n612), .B(n639), .O(n401));
  andx g381(.A(n61), .B(n675), .O(n402));
  orx  g382(.A(n411), .B(n404), .O(n403));
  orx  g383(.A(n408), .B(n405), .O(n404));
  orx  g384(.A(n407), .B(n406), .O(n405));
  andx g385(.A(n60), .B(n680), .O(n406));
  andx g386(.A(n61), .B(n669), .O(n407));
  orx  g387(.A(n410), .B(n409), .O(n408));
  andx g388(.A(n60), .B(n691), .O(n409));
  andx g389(.A(n61), .B(n43), .O(n410));
  orx  g390(.A(n418), .B(n412), .O(n411));
  orx  g391(.A(n414), .B(n413), .O(n412));
  andx g392(.A(n60), .B(n697), .O(n413));
  andx g393(.A(n61), .B(n640), .O(n414));
  orx  g394(.A(n515), .B(n416), .O(n415));
  orx  g395(.A(n455), .B(n417), .O(n416));
  orx  g396(.A(n628), .B(n508), .O(n417));
  orx  g397(.A(n481), .B(n419), .O(n418));
  andx g398(.A(n420), .B(n666), .O(n419));
  orx  g399(.A(n506), .B(n34), .O(n420));
  orx  g400(.A(n459), .B(n422), .O(po01));
  orx  g401(.A(n448), .B(n423), .O(n422));
  orx  g402(.A(n429), .B(n424), .O(n423));
  orx  g403(.A(n425), .B(n489), .O(n424));
  orx  g404(.A(n428), .B(n426), .O(n425));
  orx  g405(.A(n549), .B(n427), .O(n426));
  andx g406(.A(n21), .B(n23), .O(n427));
  andx g407(.A(n56), .B(n598), .O(n428));
  orx  g408(.A(n445), .B(n430), .O(n429));
  orx  g409(.A(n436), .B(n431), .O(n430));
  orx  g410(.A(n435), .B(n432), .O(n431));
  orx  g411(.A(n434), .B(n433), .O(n432));
  andx g412(.A(n632), .B(n53), .O(n433));
  andx g413(.A(n30), .B(n54), .O(n434));
  andx g414(.A(n33), .B(n675), .O(n435));
  orx  g415(.A(n441), .B(n437), .O(n436));
  orx  g416(.A(n440), .B(n438), .O(n437));
  andx g417(.A(n49), .B(n439), .O(n438));
  orx  g418(.A(n604), .B(n550), .O(n439));
  andx g419(.A(n598), .B(n644), .O(n440));
  orx  g420(.A(n533), .B(n442), .O(n441));
  andx g421(.A(n575), .B(n443), .O(n442));
  andx g422(.A(n444), .B(n675), .O(n443));
  orx  g423(.A(n45), .B(n631), .O(n444));
  orx  g424(.A(n447), .B(n446), .O(n445));
  andx g425(.A(n55), .B(n644), .O(n446));
  andx g426(.A(n574), .B(n604), .O(n447));
  orx  g427(.A(n452), .B(n449), .O(n448));
  orx  g428(.A(n451), .B(n450), .O(n449));
  andx g429(.A(n677), .B(n24), .O(n450));
  andx g430(.A(n650), .B(n600), .O(n451));
  orx  g431(.A(n458), .B(n453), .O(n452));
  orx  g432(.A(n456), .B(n454), .O(n453));
  andx g433(.A(n455), .B(n579), .O(n454));
  andx g434(.A(n45), .B(n629), .O(n455));
  andx g435(.A(n37), .B(n457), .O(n456));
  orx  g436(.A(n599), .B(n40), .O(n457));
  andx g437(.A(n56), .B(n601), .O(n458));
  orx  g438(.A(n473), .B(n460), .O(n459));
  orx  g439(.A(n464), .B(n461), .O(n460));
  orx  g440(.A(n463), .B(n462), .O(n461));
  andx g441(.A(n40), .B(n595), .O(n462));
  andx g442(.A(n53), .B(n581), .O(n463));
  orx  g443(.A(n470), .B(n465), .O(n464));
  orx  g444(.A(n468), .B(n466), .O(n465));
  andx g445(.A(n467), .B(n639), .O(n466));
  orx  g446(.A(n626), .B(n30), .O(n467));
  andx g447(.A(n51), .B(n469), .O(n468));
  orx  g448(.A(n602), .B(n55), .O(n469));
  andx g449(.A(n23), .B(n471), .O(n470));
  orx  g450(.A(n472), .B(n665), .O(n471));
  orx  g451(.A(n36), .B(n685), .O(n472));
  orx  g452(.A(n479), .B(n474), .O(n473));
  orx  g453(.A(n477), .B(n475), .O(n474));
  andx g454(.A(n38), .B(n476), .O(n475));
  orx  g455(.A(n669), .B(n672), .O(n476));
  andx g456(.A(n478), .B(n575), .O(n477));
  andx g457(.A(n617), .B(n45), .O(n478));
  orx  g458(.A(n484), .B(n480), .O(n479));
  orx  g459(.A(n483), .B(n481), .O(n480));
  andx g460(.A(n482), .B(n51), .O(n481));
  orx  g461(.A(n39), .B(n30), .O(n482));
  andx g462(.A(n624), .B(n617), .O(n483));
  andx g463(.A(n624), .B(n666), .O(n484));
  orx  g464(.A(n582), .B(n486), .O(po00));
  orx  g465(.A(n554), .B(n487), .O(n486));
  orx  g466(.A(n535), .B(n488), .O(n487));
  orx  g467(.A(n529), .B(n489), .O(n488));
  orx  g468(.A(n509), .B(n490), .O(n489));
  orx  g469(.A(n500), .B(n491), .O(n490));
  orx  g470(.A(n499), .B(n492), .O(n491));
  orx  g471(.A(n496), .B(n493), .O(n492));
  orx  g472(.A(n495), .B(n494), .O(n493));
  andx g473(.A(n33), .B(n632), .O(n494));
  andx g474(.A(n644), .B(n50), .O(n495));
  orx  g475(.A(n498), .B(n497), .O(n496));
  andx g476(.A(n59), .B(n669), .O(n497));
  andx g477(.A(n31), .B(n604), .O(n498));
  andx g478(.A(n23), .B(n26), .O(n499));
  orx  g479(.A(n507), .B(n501), .O(n500));
  orx  g480(.A(n503), .B(n502), .O(n501));
  andx g481(.A(n39), .B(n639), .O(n502));
  andx g482(.A(n57), .B(n504), .O(n503));
  invx g483(.A(n505), .O(n504));
  andx g484(.A(n676), .B(n618), .O(n505));
  andx g485(.A(n627), .B(n588), .O(n506));
  andx g486(.A(n508), .B(n654), .O(n507));
  andx g487(.A(n661), .B(n629), .O(n508));
  orx  g488(.A(n522), .B(n510), .O(n509));
  orx  g489(.A(n518), .B(n511), .O(n510));
  orx  g490(.A(n516), .B(n512), .O(n511));
  andx g491(.A(n515), .B(n513), .O(n512));
  orx  g492(.A(n610), .B(n514), .O(n513));
  orx  g493(.A(n649), .B(n685), .O(n514));
  andx g494(.A(n588), .B(n629), .O(n515));
  andx g495(.A(n32), .B(n517), .O(n516));
  orx  g496(.A(n43), .B(n672), .O(n517));
  andx g497(.A(n50), .B(n519), .O(n518));
  orx  g498(.A(n521), .B(n520), .O(n519));
  orx  g499(.A(n697), .B(n615), .O(n520));
  orx  g500(.A(n613), .B(n691), .O(n521));
  orx  g501(.A(n527), .B(n523), .O(n522));
  orx  g502(.A(n526), .B(n524), .O(n523));
  andx g503(.A(n646), .B(n525), .O(n524));
  orx  g504(.A(n48), .B(n54), .O(n525));
  andx g505(.A(n49), .B(n675), .O(n526));
  andx g506(.A(n617), .B(n528), .O(n527));
  orx  g507(.A(n574), .B(n33), .O(n528));
  orx  g508(.A(n534), .B(n530), .O(n529));
  orx  g509(.A(n533), .B(n531), .O(n530));
  andx g510(.A(n34), .B(n532), .O(n531));
  orx  g511(.A(n43), .B(n691), .O(n532));
  andx g512(.A(n31), .B(n26), .O(n533));
  andx g513(.A(n52), .B(n31), .O(n534));
  orx  g514(.A(n548), .B(n536), .O(n535));
  orx  g515(.A(n542), .B(n537), .O(n536));
  orx  g516(.A(n541), .B(n538), .O(n537));
  orx  g517(.A(n540), .B(n539), .O(n538));
  andx g518(.A(n30), .B(n35), .O(n539));
  andx g519(.A(n53), .B(n650), .O(n540));
  andx g520(.A(n51), .B(n34), .O(n541));
  orx  g521(.A(n547), .B(n543), .O(n542));
  orx  g522(.A(n545), .B(n544), .O(n543));
  andx g523(.A(n632), .B(n49), .O(n544));
  andx g524(.A(n40), .B(n546), .O(n545));
  orx  g525(.A(n613), .B(n56), .O(n546));
  andx g526(.A(n36), .B(n58), .O(n547));
  orx  g527(.A(n551), .B(n549), .O(n548));
  andx g528(.A(n550), .B(n59), .O(n549));
  orx  g529(.A(n632), .B(n654), .O(n550));
  andx g530(.A(n617), .B(n552), .O(n551));
  orx  g531(.A(n553), .B(n24), .O(n552));
  andx g532(.A(n575), .B(n588), .O(n553));
  orx  g533(.A(n571), .B(n555), .O(n554));
  orx  g534(.A(n567), .B(n556), .O(n555));
  orx  g535(.A(n562), .B(n557), .O(n556));
  orx  g536(.A(n559), .B(n558), .O(n557));
  andx g537(.A(n632), .B(n574), .O(n558));
  andx g538(.A(n654), .B(n560), .O(n559));
  orx  g539(.A(n33), .B(n31), .O(n560));
  andx g540(.A(n661), .B(n575), .O(n561));
  orx  g541(.A(n566), .B(n563), .O(n562));
  andx g542(.A(n56), .B(n564), .O(n563));
  orx  g543(.A(n565), .B(n34), .O(n564));
  andx g544(.A(n575), .B(n45), .O(n565));
  andx g545(.A(n26), .B(n646), .O(n566));
  orx  g546(.A(n570), .B(n568), .O(n567));
  andx g547(.A(n52), .B(n24), .O(n568));
  andx g548(.A(n588), .B(n658), .O(n569));
  andx g549(.A(n38), .B(n613), .O(n570));
  orx  g550(.A(n578), .B(n572), .O(n571));
  orx  g551(.A(n577), .B(n573), .O(n572));
  andx g552(.A(n574), .B(n675), .O(n573));
  andx g553(.A(n631), .B(n575), .O(n574));
  andx g554(.A(pi7), .B(n576), .O(n575));
  andx g555(.A(n660), .B(n707), .O(n576));
  andx g556(.A(n602), .B(n581), .O(n577));
  andx g557(.A(n628), .B(n579), .O(n578));
  orx  g558(.A(n581), .B(n580), .O(n579));
  orx  g559(.A(n604), .B(n649), .O(n580));
  orx  g560(.A(n685), .B(n610), .O(n581));
  orx  g561(.A(n606), .B(n583), .O(n582));
  orx  g562(.A(n592), .B(n584), .O(n583));
  orx  g563(.A(n590), .B(n585), .O(n584));
  andx g564(.A(n587), .B(n586), .O(n585));
  orx  g565(.A(n669), .B(n37), .O(n586));
  andx g566(.A(n588), .B(n705), .O(n587));
  invx g567(.A(n589), .O(n588));
  orx  g568(.A(n710), .B(n662), .O(n589));
  andx g569(.A(n51), .B(n591), .O(n590));
  orx  g570(.A(n646), .B(n39), .O(n591));
  orx  g571(.A(n596), .B(n593), .O(n592));
  andx g572(.A(n32), .B(n594), .O(n593));
  orx  g573(.A(n666), .B(n595), .O(n594));
  orx  g574(.A(n644), .B(n28), .O(n595));
  andx g575(.A(n604), .B(n597), .O(n596));
  orx  g576(.A(n600), .B(n598), .O(n597));
  orx  g577(.A(n599), .B(n58), .O(n598));
  andx g578(.A(n631), .B(n705), .O(n599));
  orx  g579(.A(n50), .B(n601), .O(n600));
  orx  g580(.A(n53), .B(n602), .O(n601));
  andx g581(.A(n658), .B(n45), .O(n602));
  andx g582(.A(n658), .B(n631), .O(n603));
  invx g583(.A(n605), .O(n604));
  orx  g584(.A(n701), .B(n656), .O(n605));
  orx  g585(.A(n635), .B(n607), .O(n606));
  orx  g586(.A(n622), .B(n608), .O(n607));
  andx g587(.A(n34), .B(n609), .O(n608));
  orx  g588(.A(n48), .B(n610), .O(n609));
  orx  g589(.A(n615), .B(n611), .O(n610));
  orx  g590(.A(n54), .B(n612), .O(n611));
  orx  g591(.A(n613), .B(n22), .O(n612));
  andx g592(.A(pi0), .B(n614), .O(n613));
  andx g593(.A(n703), .B(n653), .O(n614));
  orx  g594(.A(n619), .B(n616), .O(n615));
  orx  g595(.A(n617), .B(n665), .O(n616));
  invx g596(.A(n618), .O(n617));
  orx  g597(.A(n701), .B(n634), .O(n618));
  orx  g598(.A(n680), .B(n640), .O(n619));
  orx  g599(.A(n687), .B(n697), .O(n620));
  andx g600(.A(n627), .B(n45), .O(n621));
  andx g601(.A(n632), .B(n623), .O(n622));
  orx  g602(.A(n628), .B(n55), .O(n623));
  orx  g603(.A(n626), .B(n32), .O(n624));
  andx g604(.A(n627), .B(n661), .O(n625));
  andx g605(.A(n627), .B(n631), .O(n626));
  andx g606(.A(n707), .B(n659), .O(n627));
  andx g607(.A(n631), .B(n629), .O(n628));
  andx g608(.A(pi6), .B(n630), .O(n629));
  andx g609(.A(n708), .B(pi5), .O(n630));
  andx g610(.A(n662), .B(pi8), .O(n631));
  invx g611(.A(n633), .O(n632));
  orx  g612(.A(n671), .B(n634), .O(n633));
  orx  g613(.A(pi3), .B(n690), .O(n634));
  orx  g614(.A(n663), .B(n636), .O(n635));
  orx  g615(.A(n647), .B(n637), .O(n636));
  andx g616(.A(n58), .B(n638), .O(n637));
  orx  g617(.A(n644), .B(n639), .O(n638));
  orx  g618(.A(n640), .B(n42), .O(n639));
  andx g619(.A(n642), .B(n641), .O(n640));
  andx g620(.A(n690), .B(pi4), .O(n641));
  andx g621(.A(n703), .B(n643), .O(n642));
  andx g622(.A(n700), .B(n696), .O(n643));
  invx g623(.A(n645), .O(n644));
  orx  g624(.A(n671), .B(n689), .O(n645));
  andx g625(.A(n661), .B(n705), .O(n646));
  andx g626(.A(n50), .B(n648), .O(n647));
  orx  g627(.A(n654), .B(n649), .O(n648));
  orx  g628(.A(n51), .B(n42), .O(n649));
  andx g629(.A(n690), .B(n652), .O(n650));
  andx g630(.A(pi0), .B(n652), .O(n651));
  andx g631(.A(n653), .B(pi1), .O(n652));
  invx g632(.A(n694), .O(n653));
  invx g633(.A(n655), .O(n654));
  orx  g634(.A(n671), .B(n656), .O(n655));
  orx  g635(.A(pi3), .B(pi0), .O(n656));
  andx g636(.A(n661), .B(n658), .O(n657));
  andx g637(.A(n659), .B(pi5), .O(n658));
  andx g638(.A(n708), .B(n660), .O(n659));
  invx g639(.A(pi6), .O(n660));
  andx g640(.A(n662), .B(n710), .O(n661));
  invx g641(.A(pi9), .O(n662));
  andx g642(.A(n39), .B(n664), .O(n663));
  orx  g643(.A(n672), .B(n665), .O(n664));
  orx  g644(.A(n669), .B(n666), .O(n665));
  invx g645(.A(n44), .O(n666));
  orx  g646(.A(n683), .B(n668), .O(n667));
  orx  g647(.A(n690), .B(n703), .O(n668));
  invx g648(.A(n670), .O(n669));
  orx  g649(.A(n671), .B(n699), .O(n670));
  orx  g650(.A(pi1), .B(n702), .O(n671));
  orx  g651(.A(n685), .B(n673), .O(n672));
  orx  g652(.A(n35), .B(n54), .O(n673));
  orx  g653(.A(n677), .B(n37), .O(n674));
  invx g654(.A(n676), .O(n675));
  orx  g655(.A(n683), .B(n693), .O(n676));
  invx g656(.A(n678), .O(n677));
  orx  g657(.A(n683), .B(n679), .O(n678));
  orx  g658(.A(pi1), .B(n690), .O(n679));
  invx g659(.A(n681), .O(n680));
  orx  g660(.A(n683), .B(n682), .O(n681));
  orx  g661(.A(pi0), .B(n703), .O(n682));
  orx  g662(.A(n696), .B(n684), .O(n683));
  orx  g663(.A(pi4), .B(pi3), .O(n684));
  orx  g664(.A(n697), .B(n686), .O(n685));
  orx  g665(.A(n691), .B(n687), .O(n686));
  invx g666(.A(n688), .O(n687));
  orx  g667(.A(n701), .B(n689), .O(n688));
  orx  g668(.A(n700), .B(n690), .O(n689));
  invx g669(.A(pi0), .O(n690));
  invx g670(.A(n692), .O(n691));
  orx  g671(.A(n694), .B(n693), .O(n692));
  orx  g672(.A(pi1), .B(pi0), .O(n693));
  orx  g673(.A(n700), .B(n695), .O(n694));
  orx  g674(.A(pi4), .B(n696), .O(n695));
  invx g675(.A(pi2), .O(n696));
  invx g676(.A(n698), .O(n697));
  orx  g677(.A(n701), .B(n699), .O(n698));
  orx  g678(.A(pi0), .B(n700), .O(n699));
  invx g679(.A(pi3), .O(n700));
  orx  g680(.A(n703), .B(n702), .O(n701));
  orx  g681(.A(pi4), .B(pi2), .O(n702));
  invx g682(.A(pi1), .O(n703));
  andx g683(.A(n45), .B(n705), .O(n704));
  andx g684(.A(pi6), .B(n706), .O(n705));
  andx g685(.A(n708), .B(n707), .O(n706));
  invx g686(.A(pi5), .O(n707));
  invx g687(.A(pi7), .O(n708));
  andx g688(.A(n710), .B(pi9), .O(n709));
  invx g689(.A(pi8), .O(n710));
endmodule


