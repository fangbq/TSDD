
module top ( .a({\a[0][7] , \a[0][6] , \a[0][5] , \a[0][4] , \a[0][3] , 
        \a[0][2] , \a[0][1] , \a[0][0] , \a[1][7] , \a[1][6] , \a[1][5] , 
        \a[1][4] , \a[1][3] , \a[1][2] , \a[1][1] , \a[1][0] , \a[2][7] , 
        \a[2][6] , \a[2][5] , \a[2][4] , \a[2][3] , \a[2][2] , \a[2][1] , 
        \a[2][0] , \a[3][7] , \a[3][6] , \a[3][5] , \a[3][4] , \a[3][3] , 
        \a[3][2] , \a[3][1] , \a[3][0] }), y );
input \a[0][4], \a[0][5], \a[1][4], \a[1][5], \a[2][4], \a[2][5], \a[3][5], \a[3][4], \a[1][3], \a[0][3], \a[2][3], \a[3][3], \a[1][7], \a[0][7], \a[3][7], \a[2][7], \a[2][6], \a[0][6], \a[1][6], \a[3][6], \a[0][2], \a[1][2], \a[2][2], \a[3][2], \a[0][1], \a[1][1], \a[2][1], \a[3][1], \a[0][0], \a[1][0], \a[2][0], \a[3][0];  
output y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7]; 
 wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226;
  orx U1 ( .A(n1), .B(n2), .O(y[7]) );
  orx U2 ( .A(n3), .B(n4), .O(y[6]) );
  invx U3 ( .A(n5), .O(n4) );
  orx U4 ( .A(n6), .B(n7), .O(n5) );
  andx U5 ( .A(n8), .B(n7), .O(n3) );
  orx U6 ( .A(n9), .B(n10), .O(y[5]) );
  invx U7 ( .A(n11), .O(n10) );
  orx U8 ( .A(n12), .B(n13), .O(n11) );
  andx U9 ( .A(n14), .B(n13), .O(n9) );
  orx U10 ( .A(n15), .B(n16), .O(y[4]) );
  andx U11 ( .A(n17), .B(n18), .O(n16) );
  invx U12 ( .A(n19), .O(n18) );
  andx U13 ( .A(n20), .B(n19), .O(n15) );
  orx U14 ( .A(n21), .B(n22), .O(y[3]) );
  invx U15 ( .A(n23), .O(n22) );
  orx U16 ( .A(n24), .B(n25), .O(n23) );
  andx U17 ( .A(n26), .B(n25), .O(n21) );
  orx U18 ( .A(n27), .B(n28), .O(y[2]) );
  invx U19 ( .A(n29), .O(n28) );
  orx U20 ( .A(n30), .B(n31), .O(n29) );
  andx U21 ( .A(n32), .B(n31), .O(n27) );
  orx U22 ( .A(n33), .B(n34), .O(y[1]) );
  invx U23 ( .A(n35), .O(n34) );
  orx U24 ( .A(n36), .B(n37), .O(n35) );
  andx U25 ( .A(n38), .B(n37), .O(n33) );
  orx U26 ( .A(n39), .B(n40), .O(y[0]) );
  andx U27 ( .A(n41), .B(n42), .O(n40) );
  invx U28 ( .A(n43), .O(n41) );
  andx U29 ( .A(n44), .B(n43), .O(n39) );
  orx U30 ( .A(n45), .B(n37), .O(n43) );
  orx U31 ( .A(n46), .B(n31), .O(n37) );
  orx U32 ( .A(n47), .B(n25), .O(n31) );
  orx U33 ( .A(n48), .B(n19), .O(n25) );
  orx U34 ( .A(n49), .B(n13), .O(n19) );
  orx U35 ( .A(n50), .B(n7), .O(n13) );
  orx U36 ( .A(n51), .B(n52), .O(n7) );
  andx U37 ( .A(n53), .B(n1), .O(n52) );
  andx U38 ( .A(n54), .B(n55), .O(n51) );
  orx U39 ( .A(n53), .B(n1), .O(n55) );
  andx U40 ( .A(n56), .B(n57), .O(n50) );
  andx U41 ( .A(n58), .B(n59), .O(n49) );
  andx U42 ( .A(n57), .B(n20), .O(n59) );
  invx U43 ( .A(n60), .O(n58) );
  orx U44 ( .A(n17), .B(n61), .O(n60) );
  andx U45 ( .A(n62), .B(n63), .O(n48) );
  andx U46 ( .A(n64), .B(n65), .O(n47) );
  andx U47 ( .A(n63), .B(n32), .O(n65) );
  andx U48 ( .A(n30), .B(n66), .O(n64) );
  andx U49 ( .A(n67), .B(n68), .O(n46) );
  andx U50 ( .A(n36), .B(n38), .O(n67) );
  andx U51 ( .A(n69), .B(n68), .O(n45) );
  andx U52 ( .A(n66), .B(n70), .O(n68) );
  andx U53 ( .A(n71), .B(n63), .O(n70) );
  invx U54 ( .A(n72), .O(n63) );
  orx U55 ( .A(n61), .B(n73), .O(n72) );
  orx U56 ( .A(n74), .B(n75), .O(n73) );
  invx U57 ( .A(n57), .O(n75) );
  andx U58 ( .A(n76), .B(n77), .O(n57) );
  andx U59 ( .A(n78), .B(n79), .O(n77) );
  orx U60 ( .A(n8), .B(n6), .O(n79) );
  invx U61 ( .A(n53), .O(n78) );
  andx U62 ( .A(n8), .B(n6), .O(n53) );
  andx U63 ( .A(n80), .B(n81), .O(n6) );
  orx U64 ( .A(n82), .B(n83), .O(n81) );
  invx U65 ( .A(n84), .O(n80) );
  andx U66 ( .A(\a[2][6] ), .B(n83), .O(n84) );
  orx U67 ( .A(n85), .B(n86), .O(n8) );
  andx U68 ( .A(\a[1][6] ), .B(n87), .O(n86) );
  invx U69 ( .A(n88), .O(n87) );
  andx U70 ( .A(\a[0][6] ), .B(n88), .O(n85) );
  orx U71 ( .A(n1), .B(n54), .O(n76) );
  invx U72 ( .A(n2), .O(n54) );
  orx U73 ( .A(\a[2][7] ), .B(\a[3][7] ), .O(n2) );
  orx U74 ( .A(\a[0][7] ), .B(\a[1][7] ), .O(n1) );
  andx U75 ( .A(n89), .B(n17), .O(n74) );
  orx U76 ( .A(n90), .B(n91), .O(n17) );
  invx U77 ( .A(n92), .O(n91) );
  orx U78 ( .A(n93), .B(n94), .O(n92) );
  andx U79 ( .A(\a[2][4] ), .B(n94), .O(n90) );
  invx U80 ( .A(n20), .O(n89) );
  orx U81 ( .A(n95), .B(n96), .O(n20) );
  andx U82 ( .A(\a[1][4] ), .B(n97), .O(n96) );
  invx U83 ( .A(n98), .O(n97) );
  andx U84 ( .A(\a[0][4] ), .B(n98), .O(n95) );
  orx U85 ( .A(n56), .B(n99), .O(n61) );
  invx U86 ( .A(n100), .O(n99) );
  orx U87 ( .A(n12), .B(n14), .O(n100) );
  andx U88 ( .A(n14), .B(n12), .O(n56) );
  andx U89 ( .A(n101), .B(n102), .O(n12) );
  orx U90 ( .A(n103), .B(n104), .O(n102) );
  invx U91 ( .A(n105), .O(n101) );
  andx U92 ( .A(\a[2][5] ), .B(n104), .O(n105) );
  orx U93 ( .A(n106), .B(n107), .O(n14) );
  invx U94 ( .A(n108), .O(n107) );
  orx U95 ( .A(n109), .B(n110), .O(n108) );
  andx U96 ( .A(\a[0][5] ), .B(n110), .O(n106) );
  orx U97 ( .A(n32), .B(n30), .O(n71) );
  andx U98 ( .A(n111), .B(n112), .O(n30) );
  orx U99 ( .A(n113), .B(n114), .O(n112) );
  invx U100 ( .A(n115), .O(n111) );
  andx U101 ( .A(\a[2][2] ), .B(n114), .O(n115) );
  orx U102 ( .A(n116), .B(n117), .O(n32) );
  andx U103 ( .A(\a[1][2] ), .B(n118), .O(n117) );
  invx U104 ( .A(n119), .O(n118) );
  andx U105 ( .A(\a[0][2] ), .B(n119), .O(n116) );
  andx U106 ( .A(n120), .B(n121), .O(n66) );
  orx U107 ( .A(n24), .B(n26), .O(n121) );
  invx U108 ( .A(n62), .O(n120) );
  andx U109 ( .A(n26), .B(n24), .O(n62) );
  andx U110 ( .A(n122), .B(n123), .O(n24) );
  orx U111 ( .A(n124), .B(n125), .O(n123) );
  invx U112 ( .A(n126), .O(n122) );
  andx U113 ( .A(\a[2][3] ), .B(n125), .O(n126) );
  orx U114 ( .A(n127), .B(n128), .O(n26) );
  invx U115 ( .A(n129), .O(n128) );
  orx U116 ( .A(n130), .B(n131), .O(n129) );
  andx U117 ( .A(\a[0][3] ), .B(n131), .O(n127) );
  andx U118 ( .A(n132), .B(n133), .O(n69) );
  orx U119 ( .A(n36), .B(n38), .O(n133) );
  orx U120 ( .A(n134), .B(n135), .O(n38) );
  andx U121 ( .A(\a[1][1] ), .B(n136), .O(n135) );
  invx U122 ( .A(n137), .O(n136) );
  andx U123 ( .A(\a[0][1] ), .B(n137), .O(n134) );
  andx U124 ( .A(n138), .B(n139), .O(n36) );
  orx U125 ( .A(n140), .B(n141), .O(n139) );
  invx U126 ( .A(n142), .O(n138) );
  andx U127 ( .A(\a[2][1] ), .B(n141), .O(n142) );
  invx U128 ( .A(n42), .O(n132) );
  andx U129 ( .A(n143), .B(n144), .O(n42) );
  orx U130 ( .A(n145), .B(\a[2][0] ), .O(n144) );
  invx U131 ( .A(n146), .O(n145) );
  orx U132 ( .A(n146), .B(\a[3][0] ), .O(n143) );
  orx U133 ( .A(n147), .B(n141), .O(n146) );
  orx U134 ( .A(n148), .B(n114), .O(n141) );
  orx U135 ( .A(n149), .B(n125), .O(n114) );
  orx U136 ( .A(n150), .B(n94), .O(n125) );
  orx U137 ( .A(n151), .B(n104), .O(n94) );
  orx U138 ( .A(n152), .B(n83), .O(n104) );
  orx U139 ( .A(n153), .B(n154), .O(n83) );
  andx U140 ( .A(\a[2][7] ), .B(n155), .O(n154) );
  andx U141 ( .A(n156), .B(n157), .O(n153) );
  orx U142 ( .A(n155), .B(\a[2][7] ), .O(n156) );
  andx U143 ( .A(n158), .B(\a[2][5] ), .O(n152) );
  andx U144 ( .A(n159), .B(n103), .O(n158) );
  andx U145 ( .A(n160), .B(n161), .O(n151) );
  andx U146 ( .A(n162), .B(n93), .O(n161) );
  andx U147 ( .A(\a[2][4] ), .B(n159), .O(n160) );
  andx U148 ( .A(n163), .B(\a[2][3] ), .O(n150) );
  andx U149 ( .A(n164), .B(n124), .O(n163) );
  andx U150 ( .A(n165), .B(n166), .O(n149) );
  andx U151 ( .A(n164), .B(n113), .O(n166) );
  andx U152 ( .A(n167), .B(\a[2][2] ), .O(n165) );
  andx U153 ( .A(n168), .B(\a[2][1] ), .O(n148) );
  andx U154 ( .A(n169), .B(n140), .O(n168) );
  andx U155 ( .A(n170), .B(\a[2][0] ), .O(n147) );
  andx U156 ( .A(n169), .B(n171), .O(n170) );
  orx U157 ( .A(\a[2][1] ), .B(n140), .O(n171) );
  invx U158 ( .A(\a[3][1] ), .O(n140) );
  andx U159 ( .A(n167), .B(n172), .O(n169) );
  andx U160 ( .A(n173), .B(n164), .O(n172) );
  andx U161 ( .A(n159), .B(n174), .O(n164) );
  andx U162 ( .A(n162), .B(n175), .O(n174) );
  orx U163 ( .A(n93), .B(\a[2][4] ), .O(n175) );
  invx U164 ( .A(\a[3][4] ), .O(n93) );
  orx U165 ( .A(\a[2][5] ), .B(n103), .O(n162) );
  invx U166 ( .A(\a[3][5] ), .O(n103) );
  andx U167 ( .A(n176), .B(n177), .O(n159) );
  andx U168 ( .A(n178), .B(n179), .O(n177) );
  orx U169 ( .A(n82), .B(\a[2][6] ), .O(n179) );
  invx U170 ( .A(n155), .O(n178) );
  andx U171 ( .A(n82), .B(\a[2][6] ), .O(n155) );
  invx U172 ( .A(\a[3][6] ), .O(n82) );
  orx U173 ( .A(n157), .B(\a[2][7] ), .O(n176) );
  invx U174 ( .A(\a[3][7] ), .O(n157) );
  orx U175 ( .A(n113), .B(\a[2][2] ), .O(n173) );
  invx U176 ( .A(\a[3][2] ), .O(n113) );
  andx U177 ( .A(n180), .B(n181), .O(n167) );
  orx U178 ( .A(n182), .B(\a[3][3] ), .O(n181) );
  invx U179 ( .A(\a[2][3] ), .O(n182) );
  orx U180 ( .A(n124), .B(\a[2][3] ), .O(n180) );
  invx U181 ( .A(\a[3][3] ), .O(n124) );
  orx U182 ( .A(n183), .B(n184), .O(n44) );
  andx U183 ( .A(\a[1][0] ), .B(n185), .O(n184) );
  invx U184 ( .A(n186), .O(n185) );
  andx U185 ( .A(\a[0][0] ), .B(n186), .O(n183) );
  orx U186 ( .A(n187), .B(n137), .O(n186) );
  orx U187 ( .A(n188), .B(n119), .O(n137) );
  orx U188 ( .A(n189), .B(n131), .O(n119) );
  orx U189 ( .A(n190), .B(n98), .O(n131) );
  orx U190 ( .A(n191), .B(n110), .O(n98) );
  orx U191 ( .A(n192), .B(n88), .O(n110) );
  orx U192 ( .A(n193), .B(n194), .O(n88) );
  andx U193 ( .A(\a[0][7] ), .B(n195), .O(n194) );
  andx U194 ( .A(n196), .B(n197), .O(n193) );
  orx U195 ( .A(n195), .B(\a[0][7] ), .O(n196) );
  andx U196 ( .A(n198), .B(\a[0][5] ), .O(n192) );
  andx U197 ( .A(n199), .B(n109), .O(n198) );
  andx U198 ( .A(n200), .B(n201), .O(n191) );
  andx U199 ( .A(n202), .B(n203), .O(n201) );
  andx U200 ( .A(\a[0][4] ), .B(n199), .O(n200) );
  andx U201 ( .A(n204), .B(\a[0][3] ), .O(n190) );
  andx U202 ( .A(n205), .B(n130), .O(n204) );
  andx U203 ( .A(n206), .B(n207), .O(n189) );
  andx U204 ( .A(n205), .B(n208), .O(n207) );
  andx U205 ( .A(n209), .B(\a[0][2] ), .O(n206) );
  andx U206 ( .A(n210), .B(\a[0][1] ), .O(n188) );
  andx U207 ( .A(n211), .B(n212), .O(n210) );
  andx U208 ( .A(n213), .B(\a[0][0] ), .O(n187) );
  andx U209 ( .A(n211), .B(n214), .O(n213) );
  orx U210 ( .A(\a[0][1] ), .B(n212), .O(n214) );
  invx U211 ( .A(\a[1][1] ), .O(n212) );
  andx U212 ( .A(n209), .B(n215), .O(n211) );
  andx U213 ( .A(n216), .B(n205), .O(n215) );
  andx U214 ( .A(n199), .B(n217), .O(n205) );
  andx U215 ( .A(n202), .B(n218), .O(n217) );
  orx U216 ( .A(n203), .B(\a[0][4] ), .O(n218) );
  invx U217 ( .A(\a[1][4] ), .O(n203) );
  orx U218 ( .A(\a[0][5] ), .B(n109), .O(n202) );
  invx U219 ( .A(\a[1][5] ), .O(n109) );
  andx U220 ( .A(n219), .B(n220), .O(n199) );
  andx U221 ( .A(n221), .B(n222), .O(n220) );
  orx U222 ( .A(n223), .B(\a[0][6] ), .O(n222) );
  invx U223 ( .A(n195), .O(n221) );
  andx U224 ( .A(n223), .B(\a[0][6] ), .O(n195) );
  invx U225 ( .A(\a[1][6] ), .O(n223) );
  orx U226 ( .A(n197), .B(\a[0][7] ), .O(n219) );
  invx U227 ( .A(\a[1][7] ), .O(n197) );
  orx U228 ( .A(n208), .B(\a[0][2] ), .O(n216) );
  invx U229 ( .A(\a[1][2] ), .O(n208) );
  andx U230 ( .A(n224), .B(n225), .O(n209) );
  orx U231 ( .A(n226), .B(\a[1][3] ), .O(n225) );
  invx U232 ( .A(\a[0][3] ), .O(n226) );
  orx U233 ( .A(n130), .B(\a[0][3] ), .O(n224) );
  invx U234 ( .A(\a[1][3] ), .O(n130) );
endmodule

