// Benchmark "top" written by ABC on Fri Feb  7 13:38:09 2014

module top ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37,
    po0, po1, po2  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37;
  output po0, po1, po2;
  wire n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
    n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
    n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
    n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
    n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
    n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
    n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
    n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
    n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
    n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
    n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
    n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
    n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
    n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
    n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
    n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
    n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
    n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
    n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
    n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
    n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
    n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
    n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
    n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
    n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
    n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
    n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
    n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
    n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437;
  invx g0000(.a(pi03), .O(n41));
  invx g0001(.a(pi05), .O(n42));
  invx g0002(.a(pi01), .O(n43));
  invx g0003(.a(pi10), .O(n44));
  andx g0004(.a(n44), .b(n43), .O(n45));
  invx g0005(.a(pi02), .O(n46));
  invx g0006(.a(pi00), .O(n47));
  andx g0007(.a(n47), .b(n46), .O(n48));
  andx g0008(.a(n48), .b(n45), .O(n49));
  andx g0009(.a(n49), .b(n42), .O(n50));
  andx g0010(.a(n50), .b(n41), .O(n51));
  invx g0011(.a(pi07), .O(n52));
  andx g0012(.a(pi09), .b(n52), .O(n53));
  andx g0013(.a(n53), .b(pi36), .O(n54));
  andx g0014(.a(n54), .b(n51), .O(n55));
  invx g0015(.a(pi33), .O(n56));
  invx g0016(.a(pi21), .O(n57));
  andx g0017(.a(n57), .b(n56), .O(n58));
  invx g0018(.a(pi22), .O(n59));
  invx g0019(.a(pi26), .O(n60));
  andx g0020(.a(n60), .b(n59), .O(n61));
  andx g0021(.a(n61), .b(n58), .O(n62));
  invx g0022(.a(pi31), .O(n63));
  invx g0023(.a(pi29), .O(n64));
  andx g0024(.a(n64), .b(n63), .O(n65));
  invx g0025(.a(pi32), .O(n66));
  invx g0026(.a(pi12), .O(n67));
  andx g0027(.a(n67), .b(n66), .O(n68));
  andx g0028(.a(n68), .b(n65), .O(n69));
  andx g0029(.a(n69), .b(n62), .O(n70));
  andx g0030(.a(n70), .b(n55), .O(n71));
  andx g0031(.a(n63), .b(n66), .O(n72));
  andx g0032(.a(pi07), .b(n64), .O(n73));
  andx g0033(.a(n73), .b(n72), .O(n74));
  invx g0034(.a(pi06), .O(n75));
  andx g0035(.a(n59), .b(n57), .O(n76));
  andx g0036(.a(pi26), .b(n56), .O(n77));
  andx g0037(.a(n77), .b(pi10), .O(n78));
  andx g0038(.a(n78), .b(n76), .O(n79));
  invx g0039(.a(pi25), .O(n80));
  andx g0040(.a(pi17), .b(pi11), .O(n81));
  andx g0041(.a(n81), .b(n80), .O(n82));
  andx g0042(.a(n82), .b(n79), .O(n83));
  andx g0043(.a(n83), .b(n75), .O(n84));
  andx g0044(.a(n84), .b(n74), .O(n85));
  orx  g0045(.a(n85), .b(n71), .O(n86));
  invx g0046(.a(pi04), .O(n87));
  invx g0047(.a(pi20), .O(n88));
  andx g0048(.a(n80), .b(n88), .O(n89));
  andx g0049(.a(n59), .b(n66), .O(n90));
  invx g0050(.a(pi08), .O(n91));
  andx g0051(.a(n44), .b(n91), .O(n92));
  invx g0052(.a(pi13), .O(n93));
  andx g0053(.a(n93), .b(n56), .O(n94));
  andx g0054(.a(n94), .b(n92), .O(n95));
  andx g0055(.a(n95), .b(n90), .O(n96));
  andx g0056(.a(n96), .b(n89), .O(n97));
  andx g0057(.a(n97), .b(n87), .O(n98));
  invx g0058(.a(pi28), .O(n99));
  andx g0059(.a(n75), .b(n99), .O(n100));
  andx g0060(.a(pi36), .b(n63), .O(n101));
  andx g0061(.a(n101), .b(n100), .O(n102));
  andx g0062(.a(n102), .b(n98), .O(n103));
  andx g0063(.a(n59), .b(n63), .O(n104));
  andx g0064(.a(n104), .b(n66), .O(n105));
  andx g0065(.a(n105), .b(n73), .O(n106));
  invx g0066(.a(pi16), .O(n107));
  andx g0067(.a(n58), .b(n107), .O(n108));
  andx g0068(.a(n1220), .b(pi10), .O(n109));
  andx g0069(.a(n75), .b(pi11), .O(n110));
  andx g0070(.a(n110), .b(n109), .O(n111));
  andx g0071(.a(n111), .b(n106), .O(n112));
  orx  g0072(.a(n112), .b(n103), .O(n113));
  orx  g0073(.a(n113), .b(n86), .O(n114));
  andx g0074(.a(n50), .b(pi36), .O(n115));
  andx g0075(.a(n115), .b(n75), .O(n116));
  andx g0076(.a(n59), .b(n56), .O(n117));
  andx g0077(.a(n117), .b(n93), .O(n118));
  andx g0078(.a(n60), .b(n66), .O(n119));
  andx g0079(.a(n88), .b(n87), .O(n120));
  andx g0080(.a(n120), .b(n119), .O(n121));
  andx g0081(.a(n121), .b(n65), .O(n122));
  andx g0082(.a(n122), .b(n118), .O(n123));
  andx g0083(.a(n123), .b(n116), .O(n124));
  andx g0084(.a(pi07), .b(pi28), .O(n125));
  andx g0085(.a(n125), .b(n72), .O(n126));
  andx g0086(.a(n107), .b(n56), .O(n127));
  andx g0087(.a(n127), .b(pi10), .O(n128));
  andx g0088(.a(n128), .b(n76), .O(n129));
  andx g0089(.a(n80), .b(pi11), .O(n130));
  andx g0090(.a(n130), .b(n129), .O(n131));
  andx g0091(.a(n131), .b(n75), .O(n132));
  andx g0092(.a(n132), .b(n126), .O(n133));
  orx  g0093(.a(n133), .b(n124), .O(n134));
  andx g0094(.a(n51), .b(n64), .O(n135));
  andx g0095(.a(n93), .b(n57), .O(n136));
  andx g0096(.a(n136), .b(n117), .O(n137));
  andx g0097(.a(pi36), .b(n75), .O(n138));
  andx g0098(.a(n60), .b(n87), .O(n139));
  andx g0099(.a(n139), .b(n138), .O(n140));
  andx g0100(.a(n140), .b(n72), .O(n141));
  andx g0101(.a(n141), .b(n137), .O(n142));
  andx g0102(.a(n142), .b(n135), .O(n143));
  andx g0103(.a(n60), .b(n56), .O(n144));
  andx g0104(.a(n144), .b(n90), .O(n145));
  andx g0105(.a(n145), .b(pi10), .O(n146));
  andx g0106(.a(n88), .b(pi11), .O(n147));
  andx g0107(.a(n147), .b(n146), .O(n148));
  andx g0108(.a(pi17), .b(n75), .O(n149));
  andx g0109(.a(n149), .b(n148), .O(n150));
  invx g0110(.a(pi15), .O(n151));
  andx g0111(.a(pi28), .b(n151), .O(n152));
  andx g0112(.a(pi14), .b(pi07), .O(n153));
  andx g0113(.a(n153), .b(n63), .O(n154));
  andx g0114(.a(n154), .b(n152), .O(n155));
  andx g0115(.a(n155), .b(n150), .O(n156));
  orx  g0116(.a(n156), .b(n143), .O(n157));
  orx  g0117(.a(n157), .b(n134), .O(n158));
  orx  g0118(.a(n158), .b(n114), .O(n159));
  andx g0119(.a(n50), .b(n75), .O(n160));
  andx g0120(.a(n120), .b(n80), .O(n161));
  andx g0121(.a(n161), .b(n160), .O(n162));
  andx g0122(.a(n90), .b(n56), .O(n163));
  andx g0123(.a(n67), .b(n64), .O(n164));
  andx g0124(.a(n164), .b(n101), .O(n165));
  andx g0125(.a(n165), .b(n163), .O(n166));
  andx g0126(.a(n166), .b(n162), .O(n167));
  andx g0127(.a(n62), .b(pi10), .O(n168));
  andx g0128(.a(n168), .b(n81), .O(n169));
  andx g0129(.a(n169), .b(n151), .O(n170));
  andx g0130(.a(n75), .b(n66), .O(n171));
  andx g0131(.a(n171), .b(n153), .O(n172));
  andx g0132(.a(n172), .b(n65), .O(n173));
  andx g0133(.a(n173), .b(n170), .O(n174));
  orx  g0134(.a(n174), .b(n167), .O(n175));
  andx g0135(.a(n60), .b(n107), .O(n176));
  andx g0136(.a(n176), .b(pi10), .O(n177));
  andx g0137(.a(n177), .b(n117), .O(n178));
  andx g0138(.a(n178), .b(n147), .O(n179));
  andx g0139(.a(n179), .b(n75), .O(n180));
  andx g0140(.a(n180), .b(n126), .O(n181));
  andx g0141(.a(n75), .b(pi07), .O(n182));
  andx g0142(.a(n182), .b(n119), .O(n183));
  andx g0143(.a(n183), .b(n101), .O(n184));
  andx g0144(.a(n184), .b(n137), .O(n185));
  andx g0145(.a(n185), .b(n135), .O(n186));
  orx  g0146(.a(n186), .b(n181), .O(n187));
  orx  g0147(.a(n187), .b(n175), .O(n188));
  andx g0148(.a(n117), .b(n72), .O(n189));
  andx g0149(.a(n189), .b(n60), .O(n190));
  andx g0150(.a(n190), .b(pi24), .O(n191));
  andx g0151(.a(n191), .b(n88), .O(n192));
  andx g0152(.a(pi25), .b(n75), .O(n193));
  andx g0153(.a(n193), .b(n125), .O(n194));
  andx g0154(.a(n194), .b(n192), .O(n195));
  andx g0155(.a(n429), .b(n60), .O(n196));
  andx g0156(.a(n196), .b(pi27), .O(n197));
  andx g0157(.a(n99), .b(pi29), .O(n198));
  andx g0158(.a(pi09), .b(n63), .O(n199));
  andx g0159(.a(n199), .b(n52), .O(n200));
  andx g0160(.a(n200), .b(n198), .O(n201));
  andx g0161(.a(n201), .b(n197), .O(n202));
  orx  g0162(.a(n202), .b(n195), .O(n203));
  andx g0163(.a(n80), .b(n66), .O(n204));
  andx g0164(.a(n204), .b(n93), .O(n205));
  andx g0165(.a(pi07), .b(n59), .O(n206));
  andx g0166(.a(n88), .b(n56), .O(n207));
  andx g0167(.a(n207), .b(n65), .O(n208));
  andx g0168(.a(n208), .b(n206), .O(n209));
  andx g0169(.a(n209), .b(n205), .O(n210));
  andx g0170(.a(n210), .b(n116), .O(n211));
  invx g0171(.a(pi19), .O(n212));
  andx g0172(.a(n212), .b(n56), .O(n213));
  invx g0173(.a(pi18), .O(n214));
  andx g0174(.a(n60), .b(n214), .O(n215));
  andx g0175(.a(n215), .b(pi10), .O(n216));
  andx g0176(.a(n216), .b(n213), .O(n217));
  andx g0177(.a(n217), .b(n147), .O(n218));
  andx g0178(.a(n218), .b(n149), .O(n219));
  andx g0179(.a(pi28), .b(n63), .O(n220));
  andx g0180(.a(n206), .b(n66), .O(n221));
  andx g0181(.a(n221), .b(n220), .O(n222));
  andx g0182(.a(n222), .b(n219), .O(n223));
  orx  g0183(.a(n223), .b(n211), .O(n224));
  orx  g0184(.a(n224), .b(n203), .O(n225));
  orx  g0185(.a(n225), .b(n188), .O(n226));
  orx  g0186(.a(n226), .b(n159), .O(n227));
  andx g0187(.a(pi29), .b(n66), .O(n228));
  andx g0188(.a(n75), .b(n63), .O(n229));
  andx g0189(.a(n229), .b(n87), .O(n230));
  andx g0190(.a(n230), .b(n228), .O(n231));
  andx g0191(.a(n59), .b(pi30), .O(n232));
  andx g0192(.a(n232), .b(n58), .O(n233));
  andx g0193(.a(n233), .b(n60), .O(n234));
  andx g0194(.a(n234), .b(n231), .O(n235));
  andx g0195(.a(pi24), .b(n64), .O(n236));
  andx g0196(.a(n236), .b(n66), .O(n237));
  andx g0197(.a(n80), .b(n52), .O(n238));
  andx g0198(.a(n238), .b(n207), .O(n239));
  andx g0199(.a(pi23), .b(n59), .O(n240));
  andx g0200(.a(n240), .b(n199), .O(n241));
  andx g0201(.a(n241), .b(n239), .O(n242));
  andx g0202(.a(n242), .b(n237), .O(n243));
  orx  g0203(.a(n243), .b(n235), .O(n244));
  andx g0204(.a(n67), .b(pi28), .O(n245));
  andx g0205(.a(n104), .b(pi07), .O(n246));
  andx g0206(.a(n246), .b(n245), .O(n247));
  andx g0207(.a(pi23), .b(pi24), .O(n248));
  invx g0208(.a(pi11), .O(n249));
  andx g0209(.a(n249), .b(n91), .O(n250));
  andx g0210(.a(n250), .b(n75), .O(n251));
  andx g0211(.a(n251), .b(n248), .O(n252));
  andx g0212(.a(n252), .b(n247), .O(n253));
  andx g0213(.a(n75), .b(n59), .O(n254));
  andx g0214(.a(n89), .b(n56), .O(n255));
  andx g0215(.a(n255), .b(n254), .O(n256));
  andx g0216(.a(pi07), .b(pi24), .O(n257));
  andx g0217(.a(pi23), .b(n64), .O(n258));
  andx g0218(.a(n258), .b(n257), .O(n259));
  andx g0219(.a(n259), .b(n72), .O(n260));
  andx g0220(.a(n260), .b(n256), .O(n261));
  orx  g0221(.a(n261), .b(n253), .O(n262));
  orx  g0222(.a(n262), .b(n244), .O(n263));
  andx g0223(.a(n75), .b(n67), .O(n264));
  andx g0224(.a(n249), .b(pi27), .O(n265));
  andx g0225(.a(n265), .b(n264), .O(n266));
  andx g0226(.a(n99), .b(n87), .O(n267));
  andx g0227(.a(pi29), .b(n63), .O(n268));
  andx g0228(.a(n52), .b(n91), .O(n269));
  andx g0229(.a(n269), .b(n268), .O(n270));
  andx g0230(.a(n270), .b(n267), .O(n271));
  andx g0231(.a(n271), .b(n266), .O(n272));
  andx g0232(.a(n80), .b(pi29), .O(n273));
  andx g0233(.a(pi05), .b(n87), .O(n274));
  andx g0234(.a(n274), .b(n90), .O(n275));
  andx g0235(.a(n275), .b(n273), .O(n276));
  invx g0236(.a(pi27), .O(n277));
  andx g0237(.a(n277), .b(n56), .O(n278));
  andx g0238(.a(n278), .b(n88), .O(n279));
  andx g0239(.a(n229), .b(n99), .O(n280));
  andx g0240(.a(n280), .b(n279), .O(n281));
  andx g0241(.a(n281), .b(n276), .O(n282));
  orx  g0242(.a(n282), .b(n272), .O(n283));
  andx g0243(.a(n255), .b(n232), .O(n284));
  andx g0244(.a(pi07), .b(pi29), .O(n285));
  andx g0245(.a(n229), .b(n66), .O(n286));
  andx g0246(.a(n286), .b(n285), .O(n287));
  andx g0247(.a(n287), .b(n284), .O(n288));
  andx g0248(.a(n80), .b(pi28), .O(n289));
  andx g0249(.a(n289), .b(pi07), .O(n290));
  andx g0250(.a(n248), .b(n207), .O(n291));
  andx g0251(.a(n229), .b(n90), .O(n292));
  andx g0252(.a(n292), .b(n291), .O(n293));
  andx g0253(.a(n293), .b(n290), .O(n294));
  orx  g0254(.a(n294), .b(n288), .O(n295));
  orx  g0255(.a(n295), .b(n283), .O(n296));
  orx  g0256(.a(n296), .b(n263), .O(n297));
  andx g0257(.a(n93), .b(n43), .O(n298));
  andx g0258(.a(n298), .b(n48), .O(n299));
  andx g0259(.a(n299), .b(n42), .O(n300));
  andx g0260(.a(n41), .b(n249), .O(n301));
  andx g0261(.a(n301), .b(n300), .O(n302));
  invx g0262(.a(pi09), .O(n303));
  andx g0263(.a(pi36), .b(n303), .O(n304));
  andx g0264(.a(n304), .b(n75), .O(n305));
  andx g0265(.a(n305), .b(n302), .O(n306));
  andx g0266(.a(pi07), .b(n56), .O(n307));
  andx g0267(.a(n307), .b(n76), .O(n308));
  andx g0268(.a(n204), .b(n65), .O(n309));
  andx g0269(.a(n309), .b(n308), .O(n310));
  andx g0270(.a(n310), .b(n306), .O(n311));
  andx g0271(.a(n120), .b(n75), .O(n312));
  andx g0272(.a(n93), .b(n44), .O(n313));
  andx g0273(.a(n313), .b(n60), .O(n314));
  andx g0274(.a(n314), .b(n117), .O(n315));
  andx g0275(.a(n315), .b(n91), .O(n316));
  andx g0276(.a(n316), .b(n312), .O(n317));
  andx g0277(.a(pi36), .b(n66), .O(n318));
  andx g0278(.a(n318), .b(n65), .O(n319));
  andx g0279(.a(n319), .b(n317), .O(n320));
  orx  g0280(.a(n320), .b(n311), .O(n321));
  orx  g0281(.a(n321), .b(n297), .O(n322));
  andx g0282(.a(n63), .b(n56), .O(n323));
  andx g0283(.a(n323), .b(n100), .O(n324));
  andx g0284(.a(n324), .b(n76), .O(n325));
  andx g0285(.a(n44), .b(pi36), .O(n326));
  andx g0286(.a(n326), .b(n68), .O(n327));
  andx g0287(.a(n80), .b(n91), .O(n328));
  andx g0288(.a(n42), .b(n87), .O(n329));
  andx g0289(.a(n329), .b(n328), .O(n330));
  andx g0290(.a(n330), .b(n327), .O(n331));
  andx g0291(.a(n331), .b(n325), .O(n332));
  invx g0292(.a(pi30), .O(n333));
  andx g0293(.a(n333), .b(n87), .O(n334));
  andx g0294(.a(n334), .b(n171), .O(n335));
  andx g0295(.a(n207), .b(n104), .O(n336));
  andx g0296(.a(n99), .b(pi27), .O(n337));
  andx g0297(.a(n337), .b(n273), .O(n338));
  andx g0298(.a(n338), .b(n336), .O(n339));
  andx g0299(.a(n339), .b(n335), .O(n340));
  orx  g0300(.a(n340), .b(n332), .O(n341));
  andx g0301(.a(n145), .b(n92), .O(n342));
  andx g0302(.a(pi36), .b(pi07), .O(n343));
  andx g0303(.a(n343), .b(n63), .O(n344));
  andx g0304(.a(n88), .b(n64), .O(n345));
  andx g0305(.a(n345), .b(n264), .O(n346));
  andx g0306(.a(n346), .b(n344), .O(n347));
  andx g0307(.a(n347), .b(n342), .O(n348));
  andx g0308(.a(n268), .b(n59), .O(n349));
  andx g0309(.a(pi30), .b(n249), .O(n350));
  andx g0310(.a(pi07), .b(n91), .O(n351));
  andx g0311(.a(n351), .b(n350), .O(n352));
  andx g0312(.a(n352), .b(n264), .O(n353));
  andx g0313(.a(n353), .b(n349), .O(n354));
  orx  g0314(.a(n354), .b(n348), .O(n355));
  orx  g0315(.a(n355), .b(n341), .O(n356));
  andx g0316(.a(n249), .b(n64), .O(n357));
  andx g0317(.a(pi36), .b(n67), .O(n358));
  andx g0318(.a(n358), .b(n92), .O(n359));
  andx g0319(.a(n359), .b(n357), .O(n360));
  andx g0320(.a(n360), .b(n200), .O(n361));
  andx g0321(.a(n284), .b(n231), .O(n362));
  orx  g0322(.a(n362), .b(n361), .O(n363));
  andx g0323(.a(n59), .b(n67), .O(n364));
  andx g0324(.a(n364), .b(n250), .O(n365));
  andx g0325(.a(n248), .b(n182), .O(n366));
  andx g0326(.a(n366), .b(n65), .O(n367));
  andx g0327(.a(n367), .b(n365), .O(n368));
  andx g0328(.a(n60), .b(pi29), .O(n369));
  andx g0329(.a(n369), .b(n275), .O(n370));
  andx g0330(.a(n370), .b(n281), .O(n371));
  orx  g0331(.a(n371), .b(n368), .O(n372));
  orx  g0332(.a(n372), .b(n363), .O(n373));
  orx  g0333(.a(n373), .b(n356), .O(n374));
  andx g0334(.a(n144), .b(n88), .O(n375));
  andx g0335(.a(n375), .b(n232), .O(n376));
  andx g0336(.a(n376), .b(n287), .O(n377));
  andx g0337(.a(n250), .b(n63), .O(n378));
  andx g0338(.a(n378), .b(n64), .O(n379));
  andx g0339(.a(pi25), .b(n52), .O(n380));
  andx g0340(.a(pi09), .b(n67), .O(n381));
  andx g0341(.a(n381), .b(pi24), .O(n382));
  andx g0342(.a(n382), .b(n380), .O(n383));
  andx g0343(.a(n383), .b(n379), .O(n384));
  orx  g0344(.a(n384), .b(n377), .O(n385));
  andx g0345(.a(n233), .b(n80), .O(n386));
  andx g0346(.a(n386), .b(n287), .O(n387));
  andx g0347(.a(n200), .b(n228), .O(n388));
  andx g0348(.a(n388), .b(n376), .O(n389));
  orx  g0349(.a(n389), .b(n387), .O(n390));
  orx  g0350(.a(n390), .b(n385), .O(n391));
  andx g0351(.a(n238), .b(pi09), .O(n392));
  andx g0352(.a(n220), .b(n90), .O(n393));
  andx g0353(.a(n393), .b(n291), .O(n394));
  andx g0354(.a(n394), .b(n392), .O(n395));
  andx g0355(.a(n137), .b(n92), .O(n396));
  andx g0356(.a(n80), .b(n63), .O(n397));
  andx g0357(.a(n397), .b(n138), .O(n398));
  andx g0358(.a(n73), .b(n66), .O(n399));
  andx g0359(.a(n399), .b(n398), .O(n400));
  andx g0360(.a(n400), .b(n396), .O(n401));
  orx  g0361(.a(n401), .b(n395), .O(n402));
  andx g0362(.a(n337), .b(n58), .O(n403));
  andx g0363(.a(n75), .b(pi29), .O(n404));
  andx g0364(.a(n404), .b(n334), .O(n405));
  andx g0365(.a(n119), .b(n104), .O(n406));
  andx g0366(.a(n406), .b(n405), .O(n407));
  andx g0367(.a(n407), .b(n403), .O(n408));
  andx g0368(.a(n265), .b(n99), .O(n409));
  andx g0369(.a(n381), .b(n270), .O(n410));
  andx g0370(.a(n410), .b(n409), .O(n411));
  orx  g0371(.a(n411), .b(n408), .O(n412));
  orx  g0372(.a(n412), .b(n402), .O(n413));
  orx  g0373(.a(n413), .b(n391), .O(n414));
  orx  g0374(.a(n414), .b(n374), .O(n415));
  orx  g0375(.a(n415), .b(n322), .O(n416));
  andx g0376(.a(n160), .b(n80), .O(n417));
  andx g0377(.a(n318), .b(n206), .O(n418));
  andx g0378(.a(n323), .b(n164), .O(n419));
  andx g0379(.a(n419), .b(n418), .O(n420));
  andx g0380(.a(pi26), .b(n57), .O(n421));
  andx g0381(.a(n421), .b(n107), .O(n422));
  andx g0382(.a(n422), .b(n420), .O(n423));
  andx g0383(.a(n423), .b(n417), .O(n424));
  andx g0384(.a(n132), .b(n74), .O(n425));
  orx  g0385(.a(n425), .b(n424), .O(n426));
  andx g0386(.a(n302), .b(pi36), .O(n427));
  andx g0387(.a(n66), .b(n56), .O(n428));
  andx g0388(.a(n428), .b(n76), .O(n429));
  andx g0389(.a(n303), .b(n64), .O(n430));
  andx g0390(.a(n63), .b(n87), .O(n431));
  andx g0391(.a(n80), .b(n75), .O(n432));
  andx g0392(.a(n432), .b(n431), .O(n433));
  andx g0393(.a(n433), .b(n430), .O(n434));
  andx g0394(.a(n434), .b(n429), .O(n435));
  andx g0395(.a(n435), .b(n427), .O(n436));
  andx g0396(.a(n52), .b(n63), .O(n437));
  andx g0397(.a(pi36), .b(pi09), .O(n438));
  andx g0398(.a(n438), .b(n119), .O(n439));
  andx g0399(.a(n439), .b(n437), .O(n440));
  andx g0400(.a(n440), .b(n137), .O(n441));
  andx g0401(.a(n441), .b(n135), .O(n442));
  orx  g0402(.a(n442), .b(n436), .O(n443));
  orx  g0403(.a(n443), .b(n426), .O(n444));
  andx g0404(.a(n93), .b(n59), .O(n445));
  andx g0405(.a(n137), .b(n309), .O(n446));
  andx g0406(.a(n446), .b(n55), .O(n447));
  andx g0407(.a(n51), .b(pi36), .O(n448));
  andx g0408(.a(n75), .b(n64), .O(n449));
  andx g0409(.a(n431), .b(n204), .O(n450));
  andx g0410(.a(n450), .b(n449), .O(n451));
  andx g0411(.a(n451), .b(n137), .O(n452));
  andx g0412(.a(n452), .b(n448), .O(n453));
  orx  g0413(.a(n453), .b(n447), .O(n454));
  andx g0414(.a(n119), .b(n100), .O(n455));
  andx g0415(.a(n455), .b(n431), .O(n456));
  andx g0416(.a(n456), .b(n137), .O(n457));
  andx g0417(.a(n457), .b(n448), .O(n458));
  andx g0418(.a(n66), .b(n87), .O(n459));
  andx g0419(.a(n459), .b(n65), .O(n460));
  andx g0420(.a(n460), .b(n62), .O(n461));
  andx g0421(.a(n461), .b(n306), .O(n462));
  orx  g0422(.a(n462), .b(n458), .O(n463));
  orx  g0423(.a(n463), .b(n454), .O(n464));
  orx  g0424(.a(n464), .b(n444), .O(n465));
  orx  g0425(.a(n465), .b(n416), .O(n466));
  orx  g0426(.a(n466), .b(n227), .O(n467));
  andx g0427(.a(n438), .b(n50), .O(n468));
  andx g0428(.a(n468), .b(n67), .O(n469));
  andx g0429(.a(n119), .b(n107), .O(n470));
  andx g0430(.a(n214), .b(n52), .O(n471));
  andx g0431(.a(n471), .b(n76), .O(n472));
  andx g0432(.a(n213), .b(n65), .O(n473));
  andx g0433(.a(n473), .b(n472), .O(n474));
  andx g0434(.a(n474), .b(n470), .O(n475));
  andx g0435(.a(n475), .b(n469), .O(n476));
  andx g0436(.a(n343), .b(n51), .O(n477));
  andx g0437(.a(n76), .b(n93), .O(n478));
  andx g0438(.a(n428), .b(n397), .O(n479));
  andx g0439(.a(n479), .b(n449), .O(n480));
  andx g0440(.a(n480), .b(n478), .O(n481));
  andx g0441(.a(n481), .b(n477), .O(n482));
  orx  g0442(.a(n482), .b(n476), .O(n483));
  andx g0443(.a(n88), .b(n93), .O(n484));
  andx g0444(.a(n328), .b(n249), .O(n485));
  andx g0445(.a(n485), .b(n484), .O(n486));
  andx g0446(.a(n486), .b(n189), .O(n487));
  andx g0447(.a(n487), .b(n87), .O(n488));
  andx g0448(.a(n430), .b(n138), .O(n489));
  andx g0449(.a(n489), .b(n488), .O(n490));
  andx g0450(.a(n80), .b(n87), .O(n491));
  andx g0451(.a(n491), .b(n100), .O(n492));
  andx g0452(.a(n492), .b(n51), .O(n493));
  andx g0453(.a(n57), .b(n66), .O(n494));
  andx g0454(.a(n494), .b(n56), .O(n495));
  andx g0455(.a(n364), .b(n101), .O(n496));
  andx g0456(.a(n496), .b(n495), .O(n497));
  andx g0457(.a(n497), .b(n493), .O(n498));
  orx  g0458(.a(n498), .b(n490), .O(n499));
  orx  g0459(.a(n499), .b(n483), .O(n500));
  andx g0460(.a(n196), .b(pi24), .O(n501));
  andx g0461(.a(n431), .b(n193), .O(n502));
  andx g0462(.a(n502), .b(n501), .O(n503));
  andx g0463(.a(n51), .b(n67), .O(n504));
  andx g0464(.a(n138), .b(n65), .O(n505));
  andx g0465(.a(n505), .b(n491), .O(n506));
  andx g0466(.a(n506), .b(n429), .O(n507));
  andx g0467(.a(n507), .b(n504), .O(n508));
  orx  g0468(.a(n508), .b(n503), .O(n509));
  andx g0469(.a(n52), .b(n59), .O(n510));
  andx g0470(.a(n510), .b(n119), .O(n511));
  andx g0471(.a(n511), .b(n208), .O(n512));
  andx g0472(.a(n512), .b(n469), .O(n513));
  andx g0473(.a(pi36), .b(n99), .O(n514));
  andx g0474(.a(n514), .b(n72), .O(n515));
  andx g0475(.a(n515), .b(n317), .O(n516));
  orx  g0476(.a(n516), .b(n513), .O(n517));
  orx  g0477(.a(n517), .b(n509), .O(n518));
  orx  g0478(.a(n518), .b(n500), .O(n519));
  andx g0479(.a(n50), .b(n67), .O(n520));
  andx g0480(.a(n520), .b(n75), .O(n521));
  andx g0481(.a(n65), .b(pi07), .O(n522));
  andx g0482(.a(n80), .b(pi36), .O(n523));
  andx g0483(.a(n207), .b(n90), .O(n524));
  andx g0484(.a(n524), .b(n523), .O(n525));
  andx g0485(.a(n525), .b(n522), .O(n526));
  andx g0486(.a(n526), .b(n521), .O(n527));
  andx g0487(.a(n304), .b(n100), .O(n528));
  andx g0488(.a(n528), .b(n488), .O(n529));
  andx g0489(.a(n126), .b(n84), .O(n530));
  orx  g0490(.a(n530), .b(n529), .O(n531));
  orx  g0491(.a(n531), .b(n527), .O(n532));
  invx g0492(.a(pi17), .O(n533));
  andx g0493(.a(n160), .b(n533), .O(n534));
  andx g0494(.a(n307), .b(n93), .O(n535));
  andx g0495(.a(n107), .b(n57), .O(n536));
  andx g0496(.a(n536), .b(n318), .O(n537));
  andx g0497(.a(n60), .b(n64), .O(n538));
  andx g0498(.a(n538), .b(n104), .O(n539));
  andx g0499(.a(n539), .b(n537), .O(n540));
  andx g0500(.a(n540), .b(n535), .O(n541));
  andx g0501(.a(n541), .b(n534), .O(n542));
  andx g0502(.a(n300), .b(n88), .O(n543));
  andx g0503(.a(n543), .b(n138), .O(n544));
  andx g0504(.a(n303), .b(pi07), .O(n545));
  andx g0505(.a(n397), .b(n357), .O(n546));
  andx g0506(.a(n546), .b(n545), .O(n547));
  andx g0507(.a(n547), .b(n163), .O(n548));
  andx g0508(.a(n548), .b(n544), .O(n549));
  orx  g0509(.a(n549), .b(n542), .O(n550));
  andx g0510(.a(n90), .b(n60), .O(n551));
  andx g0511(.a(pi36), .b(n56), .O(n552));
  andx g0512(.a(n552), .b(n65), .O(n553));
  andx g0513(.a(n553), .b(n120), .O(n554));
  andx g0514(.a(n554), .b(n551), .O(n555));
  andx g0515(.a(n555), .b(n521), .O(n556));
  andx g0516(.a(n249), .b(n87), .O(n557));
  andx g0517(.a(n557), .b(n323), .O(n558));
  andx g0518(.a(n558), .b(n430), .O(n559));
  andx g0519(.a(n559), .b(n551), .O(n560));
  andx g0520(.a(n560), .b(n544), .O(n561));
  orx  g0521(.a(n561), .b(n556), .O(n562));
  orx  g0522(.a(n562), .b(n550), .O(n563));
  orx  g0523(.a(n563), .b(n532), .O(n564));
  orx  g0524(.a(n564), .b(n519), .O(n565));
  andx g0525(.a(pi14), .b(n151), .O(n566));
  andx g0526(.a(n522), .b(n566), .O(n567));
  andx g0527(.a(n567), .b(n150), .O(n568));
  andx g0528(.a(n552), .b(n72), .O(n569));
  andx g0529(.a(n569), .b(n478), .O(n570));
  andx g0530(.a(n570), .b(n493), .O(n571));
  orx  g0531(.a(n571), .b(n568), .O(n572));
  andx g0532(.a(n60), .b(n57), .O(n573));
  andx g0533(.a(n573), .b(n107), .O(n574));
  andx g0534(.a(n574), .b(n420), .O(n575));
  andx g0535(.a(n575), .b(n534), .O(n576));
  andx g0536(.a(n76), .b(n60), .O(n577));
  andx g0537(.a(n428), .b(n229), .O(n578));
  andx g0538(.a(n578), .b(n164), .O(n579));
  andx g0539(.a(n579), .b(n577), .O(n580));
  andx g0540(.a(n580), .b(n477), .O(n581));
  orx  g0541(.a(n581), .b(n576), .O(n582));
  orx  g0542(.a(n582), .b(n572), .O(n583));
  andx g0543(.a(pi09), .b(pi28), .O(n584));
  andx g0544(.a(n584), .b(n380), .O(n585));
  andx g0545(.a(n585), .b(n192), .O(n586));
  andx g0546(.a(n115), .b(n67), .O(n587));
  andx g0547(.a(n72), .b(n56), .O(n588));
  andx g0548(.a(n59), .b(n64), .O(n589));
  andx g0549(.a(n589), .b(n89), .O(n590));
  andx g0550(.a(n590), .b(n53), .O(n591));
  andx g0551(.a(n591), .b(n588), .O(n592));
  andx g0552(.a(n592), .b(n587), .O(n593));
  orx  g0553(.a(n593), .b(n586), .O(n594));
  andx g0554(.a(n285), .b(n63), .O(n595));
  andx g0555(.a(n595), .b(n100), .O(n596));
  andx g0556(.a(n596), .b(n197), .O(n597));
  andx g0557(.a(n222), .b(n111), .O(n598));
  orx  g0558(.a(n598), .b(n597), .O(n599));
  orx  g0559(.a(n599), .b(n594), .O(n600));
  orx  g0560(.a(n600), .b(n583), .O(n601));
  andx g0561(.a(n77), .b(n93), .O(n602));
  andx g0562(.a(n104), .b(n73), .O(n603));
  andx g0563(.a(n603), .b(n537), .O(n604));
  andx g0564(.a(n604), .b(n602), .O(n605));
  andx g0565(.a(n605), .b(n417), .O(n606));
  andx g0566(.a(n219), .b(n106), .O(n607));
  orx  g0567(.a(n607), .b(n606), .O(n608));
  andx g0568(.a(pi14), .b(pi09), .O(n609));
  andx g0569(.a(pi28), .b(n66), .O(n610));
  andx g0570(.a(n610), .b(n609), .O(n611));
  andx g0571(.a(n611), .b(n437), .O(n612));
  andx g0572(.a(n612), .b(n170), .O(n613));
  andx g0573(.a(n505), .b(n98), .O(n614));
  orx  g0574(.a(n614), .b(n613), .O(n615));
  orx  g0575(.a(n615), .b(n608), .O(n616));
  andx g0576(.a(n139), .b(n58), .O(n617));
  andx g0577(.a(n303), .b(n99), .O(n618));
  andx g0578(.a(n292), .b(n618), .O(n619));
  andx g0579(.a(n619), .b(n617), .O(n620));
  andx g0580(.a(n620), .b(n427), .O(n621));
  andx g0581(.a(n180), .b(n74), .O(n622));
  orx  g0582(.a(n622), .b(n621), .O(n623));
  andx g0583(.a(n494), .b(n61), .O(n624));
  andx g0584(.a(n323), .b(n267), .O(n625));
  andx g0585(.a(n625), .b(n138), .O(n626));
  andx g0586(.a(n626), .b(n624), .O(n627));
  andx g0587(.a(n627), .b(n504), .O(n628));
  andx g0588(.a(n90), .b(n93), .O(n629));
  andx g0589(.a(n629), .b(n553), .O(n630));
  andx g0590(.a(n630), .b(n162), .O(n631));
  orx  g0591(.a(n631), .b(n628), .O(n632));
  orx  g0592(.a(n632), .b(n623), .O(n633));
  orx  g0593(.a(n633), .b(n616), .O(n634));
  orx  g0594(.a(n634), .b(n601), .O(n635));
  orx  g0595(.a(n635), .b(n565), .O(n636));
  orx  g0596(.a(n636), .b(n467), .O(n637));
  andx g0597(.a(n216), .b(n58), .O(n638));
  andx g0598(.a(n638), .b(n81), .O(n639));
  andx g0599(.a(n104), .b(n212), .O(n640));
  andx g0600(.a(n610), .b(n53), .O(n641));
  andx g0601(.a(n641), .b(n640), .O(n642));
  andx g0602(.a(n642), .b(n639), .O(n643));
  andx g0603(.a(n93), .b(n64), .O(n644));
  andx g0604(.a(n644), .b(n428), .O(n645));
  andx g0605(.a(n536), .b(n53), .O(n646));
  andx g0606(.a(n60), .b(n533), .O(n647));
  andx g0607(.a(n647), .b(n104), .O(n648));
  andx g0608(.a(n648), .b(n646), .O(n649));
  andx g0609(.a(n649), .b(n645), .O(n650));
  andx g0610(.a(n650), .b(n115), .O(n651));
  orx  g0611(.a(n651), .b(n643), .O(n652));
  andx g0612(.a(n72), .b(pi07), .O(n653));
  andx g0613(.a(n345), .b(n138), .O(n654));
  andx g0614(.a(n654), .b(n653), .O(n655));
  andx g0615(.a(n655), .b(n316), .O(n656));
  andx g0616(.a(n92), .b(n89), .O(n657));
  andx g0617(.a(n657), .b(n189), .O(n658));
  andx g0618(.a(n658), .b(n87), .O(n659));
  andx g0619(.a(pi36), .b(n64), .O(n660));
  andx g0620(.a(n660), .b(n264), .O(n661));
  andx g0621(.a(n661), .b(n659), .O(n662));
  orx  g0622(.a(n662), .b(n656), .O(n663));
  orx  g0623(.a(n663), .b(n652), .O(n664));
  andx g0624(.a(n128), .b(n90), .O(n665));
  andx g0625(.a(n147), .b(n80), .O(n666));
  andx g0626(.a(n666), .b(n665), .O(n667));
  andx g0627(.a(n65), .b(n53), .O(n668));
  andx g0628(.a(n668), .b(n667), .O(n669));
  andx g0629(.a(n220), .b(n182), .O(n670));
  andx g0630(.a(n670), .b(n667), .O(n671));
  orx  g0631(.a(n671), .b(n669), .O(n672));
  andx g0632(.a(n522), .b(n138), .O(n673));
  andx g0633(.a(n673), .b(n97), .O(n674));
  andx g0634(.a(n107), .b(n43), .O(n675));
  andx g0635(.a(n48), .b(n44), .O(n676));
  andx g0636(.a(n676), .b(n675), .O(n677));
  andx g0637(.a(n677), .b(n87), .O(n678));
  andx g0638(.a(pi29), .b(n57), .O(n679));
  andx g0639(.a(n679), .b(n61), .O(n680));
  andx g0640(.a(n533), .b(n99), .O(n681));
  andx g0641(.a(n681), .b(n101), .O(n682));
  andx g0642(.a(n428), .b(n264), .O(n683));
  andx g0643(.a(n683), .b(n682), .O(n684));
  andx g0644(.a(n684), .b(n680), .O(n685));
  andx g0645(.a(n685), .b(n678), .O(n686));
  orx  g0646(.a(n686), .b(n674), .O(n687));
  orx  g0647(.a(n687), .b(n672), .O(n688));
  orx  g0648(.a(n688), .b(n664), .O(n689));
  andx g0649(.a(n437), .b(n66), .O(n690));
  andx g0650(.a(n690), .b(n584), .O(n691));
  andx g0651(.a(n691), .b(n179), .O(n692));
  andx g0652(.a(n437), .b(n59), .O(n693));
  andx g0653(.a(pi11), .b(n66), .O(n694));
  andx g0654(.a(n694), .b(n584), .O(n695));
  andx g0655(.a(n695), .b(n693), .O(n696));
  andx g0656(.a(n696), .b(n109), .O(n697));
  orx  g0657(.a(n697), .b(n692), .O(n698));
  andx g0658(.a(n76), .b(n56), .O(n699));
  andx g0659(.a(n699), .b(n72), .O(n700));
  andx g0660(.a(n700), .b(n248), .O(n701));
  andx g0661(.a(n584), .b(n238), .O(n702));
  andx g0662(.a(n702), .b(n701), .O(n703));
  andx g0663(.a(n80), .b(pi27), .O(n704));
  andx g0664(.a(n704), .b(n700), .O(n705));
  andx g0665(.a(n285), .b(n100), .O(n706));
  andx g0666(.a(n706), .b(n705), .O(n707));
  orx  g0667(.a(n707), .b(n703), .O(n708));
  orx  g0668(.a(n708), .b(n698), .O(n709));
  andx g0669(.a(n198), .b(n53), .O(n710));
  andx g0670(.a(n710), .b(n705), .O(n711));
  andx g0671(.a(n65), .b(n59), .O(n712));
  andx g0672(.a(n694), .b(n53), .O(n713));
  andx g0673(.a(n713), .b(n712), .O(n714));
  andx g0674(.a(n714), .b(n109), .O(n715));
  orx  g0675(.a(n715), .b(n711), .O(n716));
  andx g0676(.a(n1220), .b(pi05), .O(n717));
  andx g0677(.a(n59), .b(pi29), .O(n718));
  andx g0678(.a(n718), .b(n431), .O(n719));
  andx g0679(.a(n681), .b(n171), .O(n720));
  andx g0680(.a(n720), .b(n719), .O(n721));
  andx g0681(.a(n721), .b(n717), .O(n722));
  andx g0682(.a(n432), .b(n125), .O(n723));
  andx g0683(.a(n723), .b(n701), .O(n724));
  orx  g0684(.a(n724), .b(n722), .O(n725));
  orx  g0685(.a(n725), .b(n716), .O(n726));
  orx  g0686(.a(n726), .b(n709), .O(n727));
  orx  g0687(.a(n727), .b(n689), .O(n728));
  andx g0688(.a(n48), .b(n93), .O(n729));
  andx g0689(.a(n729), .b(n675), .O(n730));
  andx g0690(.a(n100), .b(n87), .O(n731));
  andx g0691(.a(n731), .b(n730), .O(n732));
  andx g0692(.a(pi14), .b(n56), .O(n733));
  andx g0693(.a(n733), .b(n679), .O(n734));
  andx g0694(.a(n151), .b(n63), .O(n735));
  andx g0695(.a(n735), .b(n304), .O(n736));
  andx g0696(.a(n736), .b(n734), .O(n737));
  andx g0697(.a(n737), .b(n551), .O(n738));
  andx g0698(.a(n738), .b(n732), .O(n739));
  andx g0699(.a(n538), .b(n264), .O(n740));
  andx g0700(.a(n740), .b(n733), .O(n741));
  andx g0701(.a(n107), .b(n151), .O(n742));
  andx g0702(.a(n742), .b(n76), .O(n743));
  andx g0703(.a(n343), .b(n72), .O(n744));
  andx g0704(.a(n744), .b(n743), .O(n745));
  andx g0705(.a(n745), .b(n741), .O(n746));
  andx g0706(.a(n746), .b(n50), .O(n747));
  orx  g0707(.a(n747), .b(n739), .O(n748));
  andx g0708(.a(n80), .b(pi26), .O(n749));
  andx g0709(.a(n749), .b(n679), .O(n750));
  andx g0710(.a(n67), .b(n99), .O(n751));
  andx g0711(.a(n751), .b(n138), .O(n752));
  andx g0712(.a(n752), .b(n189), .O(n753));
  andx g0713(.a(n753), .b(n750), .O(n754));
  andx g0714(.a(n754), .b(n678), .O(n755));
  andx g0715(.a(n52), .b(n64), .O(n756));
  andx g0716(.a(n756), .b(n735), .O(n757));
  andx g0717(.a(n757), .b(n609), .O(n758));
  andx g0718(.a(n144), .b(n93), .O(n759));
  andx g0719(.a(n536), .b(n90), .O(n760));
  andx g0720(.a(n760), .b(n759), .O(n761));
  andx g0721(.a(n761), .b(n758), .O(n762));
  andx g0722(.a(n762), .b(n115), .O(n763));
  orx  g0723(.a(n763), .b(n755), .O(n764));
  orx  g0724(.a(n764), .b(n748), .O(n765));
  andx g0725(.a(n430), .b(pi07), .O(n766));
  andx g0726(.a(n766), .b(n138), .O(n767));
  andx g0727(.a(n767), .b(n487), .O(n768));
  andx g0728(.a(n730), .b(n87), .O(n769));
  andx g0729(.a(pi26), .b(n59), .O(n770));
  andx g0730(.a(n770), .b(n273), .O(n771));
  andx g0731(.a(n100), .b(n58), .O(n772));
  andx g0732(.a(n304), .b(n72), .O(n773));
  andx g0733(.a(n773), .b(n772), .O(n774));
  andx g0734(.a(n774), .b(n771), .O(n775));
  andx g0735(.a(n775), .b(n769), .O(n776));
  orx  g0736(.a(n776), .b(n768), .O(n777));
  andx g0737(.a(n62), .b(n93), .O(n778));
  andx g0738(.a(n778), .b(n250), .O(n779));
  andx g0739(.a(n430), .b(n66), .O(n780));
  andx g0740(.a(n431), .b(n138), .O(n781));
  andx g0741(.a(n781), .b(n780), .O(n782));
  andx g0742(.a(n782), .b(n779), .O(n783));
  andx g0743(.a(pi17), .b(n52), .O(n784));
  andx g0744(.a(n784), .b(n584), .O(n785));
  andx g0745(.a(n785), .b(n105), .O(n786));
  andx g0746(.a(n786), .b(n218), .O(n787));
  orx  g0747(.a(n787), .b(n783), .O(n788));
  orx  g0748(.a(n788), .b(n777), .O(n789));
  orx  g0749(.a(n789), .b(n765), .O(n790));
  andx g0750(.a(n691), .b(n83), .O(n791));
  andx g0751(.a(n90), .b(n78), .O(n792));
  andx g0752(.a(n80), .b(pi17), .O(n793));
  andx g0753(.a(n793), .b(n147), .O(n794));
  andx g0754(.a(n794), .b(n792), .O(n795));
  andx g0755(.a(n795), .b(n668), .O(n796));
  orx  g0756(.a(n796), .b(n791), .O(n797));
  andx g0757(.a(n438), .b(n345), .O(n798));
  andx g0758(.a(n798), .b(n690), .O(n799));
  andx g0759(.a(n799), .b(n316), .O(n800));
  andx g0760(.a(n72), .b(n212), .O(n801));
  andx g0761(.a(n254), .b(n73), .O(n802));
  andx g0762(.a(n802), .b(n801), .O(n803));
  andx g0763(.a(n803), .b(n639), .O(n804));
  orx  g0764(.a(n804), .b(n800), .O(n805));
  orx  g0765(.a(n805), .b(n797), .O(n806));
  andx g0766(.a(n536), .b(n117), .O(n807));
  andx g0767(.a(n749), .b(n438), .O(n808));
  andx g0768(.a(n756), .b(n72), .O(n809));
  andx g0769(.a(n809), .b(n808), .O(n810));
  andx g0770(.a(n810), .b(n807), .O(n811));
  andx g0771(.a(n811), .b(n520), .O(n812));
  andx g0772(.a(n675), .b(n48), .O(n813));
  andx g0773(.a(n813), .b(n42), .O(n814));
  andx g0774(.a(n814), .b(n87), .O(n815));
  andx g0775(.a(n647), .b(n494), .O(n816));
  andx g0776(.a(n264), .b(n117), .O(n817));
  andx g0777(.a(n304), .b(n65), .O(n818));
  andx g0778(.a(n818), .b(n817), .O(n819));
  andx g0779(.a(n819), .b(n816), .O(n820));
  andx g0780(.a(n820), .b(n815), .O(n821));
  orx  g0781(.a(n821), .b(n812), .O(n822));
  andx g0782(.a(n653), .b(n489), .O(n823));
  andx g0783(.a(n823), .b(n779), .O(n824));
  andx g0784(.a(n343), .b(n75), .O(n825));
  andx g0785(.a(n825), .b(n50), .O(n826));
  andx g0786(.a(n538), .b(n445), .O(n827));
  andx g0787(.a(n207), .b(n72), .O(n828));
  andx g0788(.a(n828), .b(n827), .O(n829));
  andx g0789(.a(n829), .b(n826), .O(n830));
  orx  g0790(.a(n830), .b(n824), .O(n831));
  orx  g0791(.a(n831), .b(n822), .O(n832));
  orx  g0792(.a(n832), .b(n806), .O(n833));
  orx  g0793(.a(n833), .b(n790), .O(n834));
  orx  g0794(.a(n834), .b(n728), .O(n835));
  andx g0795(.a(n448), .b(n264), .O(n836));
  andx g0796(.a(n139), .b(n72), .O(n837));
  andx g0797(.a(n461), .b(n836), .O(n838));
  andx g0798(.a(n587), .b(n75), .O(n839));
  andx g0799(.a(n214), .b(n57), .O(n840));
  andx g0800(.a(n840), .b(n213), .O(n841));
  andx g0801(.a(n603), .b(n841), .O(n842));
  andx g0802(.a(n842), .b(n470), .O(n843));
  andx g0803(.a(n843), .b(n839), .O(n844));
  andx g0804(.a(n501), .b(pi25), .O(n845));
  andx g0805(.a(n845), .b(n670), .O(n846));
  orx  g0806(.a(n846), .b(n844), .O(n847));
  orx  g0807(.a(n847), .b(n838), .O(n848));
  andx g0808(.a(n206), .b(n119), .O(n849));
  andx g0809(.a(n849), .b(n208), .O(n850));
  andx g0810(.a(n850), .b(n839), .O(n851));
  andx g0811(.a(n343), .b(n264), .O(n852));
  andx g0812(.a(n852), .b(n566), .O(n853));
  andx g0813(.a(n589), .b(n573), .O(n854));
  andx g0814(.a(n303), .b(n63), .O(n855));
  andx g0815(.a(n855), .b(n428), .O(n856));
  andx g0816(.a(n856), .b(n854), .O(n857));
  andx g0817(.a(n857), .b(n853), .O(n858));
  andx g0818(.a(n858), .b(n814), .O(n859));
  andx g0819(.a(n54), .b(n50), .O(n860));
  andx g0820(.a(n214), .b(n107), .O(n861));
  andx g0821(.a(n861), .b(n93), .O(n862));
  andx g0822(.a(n538), .b(n213), .O(n863));
  andx g0823(.a(n76), .b(n72), .O(n864));
  andx g0824(.a(n864), .b(n863), .O(n865));
  andx g0825(.a(n865), .b(n862), .O(n866));
  andx g0826(.a(n866), .b(n860), .O(n867));
  andx g0827(.a(n731), .b(n677), .O(n868));
  andx g0828(.a(n117), .b(n60), .O(n869));
  andx g0829(.a(n679), .b(n566), .O(n870));
  andx g0830(.a(n101), .b(n68), .O(n871));
  andx g0831(.a(n871), .b(n870), .O(n872));
  andx g0832(.a(n872), .b(n869), .O(n873));
  andx g0833(.a(n873), .b(n868), .O(n874));
  orx  g0834(.a(n874), .b(n867), .O(n875));
  orx  g0835(.a(n875), .b(n859), .O(n876));
  orx  g0836(.a(n876), .b(n851), .O(n877));
  andx g0837(.a(n584), .b(n437), .O(n878));
  andx g0838(.a(n878), .b(n845), .O(n879));
  andx g0839(.a(n310), .b(n836), .O(n880));
  orx  g0840(.a(n880), .b(n879), .O(n881));
  orx  g0841(.a(n881), .b(n877), .O(n882));
  orx  g0842(.a(n882), .b(n848), .O(n883));
  orx  g0843(.a(n883), .b(n835), .O(n884));
  andx g0844(.a(n647), .b(n199), .O(n885));
  andx g0845(.a(n756), .b(n318), .O(n886));
  andx g0846(.a(n886), .b(n885), .O(n887));
  andx g0847(.a(n887), .b(n807), .O(n888));
  andx g0848(.a(n888), .b(n520), .O(n889));
  andx g0849(.a(n43), .b(n56), .O(n890));
  andx g0850(.a(n890), .b(n48), .O(n891));
  andx g0851(.a(n891), .b(n42), .O(n892));
  andx g0852(.a(n892), .b(n301), .O(n893));
  andx g0853(.a(n431), .b(n57), .O(n894));
  andx g0854(.a(n303), .b(n67), .O(n895));
  andx g0855(.a(n895), .b(n204), .O(n896));
  andx g0856(.a(n514), .b(n254), .O(n897));
  andx g0857(.a(n897), .b(n896), .O(n898));
  andx g0858(.a(n898), .b(n894), .O(n899));
  andx g0859(.a(n899), .b(n893), .O(n900));
  orx  g0860(.a(n900), .b(n889), .O(n901));
  andx g0861(.a(pi09), .b(n64), .O(n902));
  andx g0862(.a(n902), .b(n63), .O(n903));
  andx g0863(.a(n784), .b(n566), .O(n904));
  andx g0864(.a(n904), .b(n903), .O(n905));
  andx g0865(.a(n905), .b(n148), .O(n906));
  andx g0866(.a(n58), .b(n44), .O(n907));
  andx g0867(.a(n907), .b(n93), .O(n908));
  andx g0868(.a(n42), .b(n59), .O(n909));
  andx g0869(.a(n909), .b(n328), .O(n910));
  andx g0870(.a(n910), .b(n459), .O(n911));
  andx g0871(.a(n911), .b(n102), .O(n912));
  andx g0872(.a(n912), .b(n908), .O(n913));
  orx  g0873(.a(n913), .b(n906), .O(n914));
  orx  g0874(.a(n914), .b(n901), .O(n915));
  andx g0875(.a(n752), .b(n659), .O(n916));
  andx g0876(.a(pi17), .b(n66), .O(n917));
  andx g0877(.a(n917), .b(n53), .O(n918));
  andx g0878(.a(n918), .b(n712), .O(n919));
  andx g0879(.a(n919), .b(n218), .O(n920));
  orx  g0880(.a(n920), .b(n916), .O(n921));
  andx g0881(.a(n48), .b(n43), .O(n922));
  andx g0882(.a(n922), .b(n861), .O(n923));
  andx g0883(.a(n459), .b(n404), .O(n924));
  andx g0884(.a(n924), .b(n751), .O(n925));
  andx g0885(.a(n60), .b(n212), .O(n926));
  andx g0886(.a(n926), .b(n76), .O(n927));
  andx g0887(.a(n855), .b(n552), .O(n928));
  andx g0888(.a(n928), .b(n927), .O(n929));
  andx g0889(.a(n929), .b(n925), .O(n930));
  andx g0890(.a(n930), .b(n923), .O(n931));
  andx g0891(.a(n431), .b(n171), .O(n932));
  andx g0892(.a(n932), .b(n304), .O(n933));
  andx g0893(.a(n215), .b(n127), .O(n934));
  andx g0894(.a(n212), .b(n57), .O(n935));
  andx g0895(.a(n935), .b(n589), .O(n936));
  andx g0896(.a(n936), .b(n934), .O(n937));
  andx g0897(.a(n937), .b(n933), .O(n938));
  andx g0898(.a(n938), .b(n300), .O(n939));
  orx  g0899(.a(n939), .b(n931), .O(n940));
  orx  g0900(.a(n940), .b(n921), .O(n941));
  orx  g0901(.a(n941), .b(n915), .O(n942));
  andx g0902(.a(n676), .b(n298), .O(n943));
  andx g0903(.a(n138), .b(n120), .O(n944));
  andx g0904(.a(n59), .b(n99), .O(n945));
  andx g0905(.a(n945), .b(n273), .O(n946));
  andx g0906(.a(n946), .b(n944), .O(n947));
  andx g0907(.a(n947), .b(n588), .O(n948));
  andx g0908(.a(n948), .b(n943), .O(n949));
  andx g0909(.a(n618), .b(n204), .O(n950));
  andx g0910(.a(n950), .b(n781), .O(n951));
  andx g0911(.a(n951), .b(n699), .O(n952));
  andx g0912(.a(n952), .b(n302), .O(n953));
  orx  g0913(.a(n953), .b(n949), .O(n954));
  andx g0914(.a(n220), .b(n212), .O(n955));
  andx g0915(.a(n206), .b(n171), .O(n956));
  andx g0916(.a(n956), .b(n955), .O(n957));
  andx g0917(.a(n957), .b(n639), .O(n958));
  andx g0918(.a(n437), .b(n204), .O(n959));
  andx g0919(.a(n902), .b(n358), .O(n960));
  andx g0920(.a(n960), .b(n959), .O(n961));
  andx g0921(.a(n961), .b(n699), .O(n962));
  andx g0922(.a(n962), .b(n51), .O(n963));
  orx  g0923(.a(n963), .b(n958), .O(n964));
  orx  g0924(.a(n964), .b(n954), .O(n965));
  andx g0925(.a(n342), .b(n312), .O(n966));
  andx g0926(.a(n165), .b(n966), .O(n967));
  andx g0927(.a(n566), .b(n489), .O(n968));
  andx g0928(.a(n837), .b(n807), .O(n969));
  andx g0929(.a(n969), .b(n968), .O(n970));
  andx g0930(.a(n970), .b(n300), .O(n971));
  orx  g0931(.a(n971), .b(n967), .O(n972));
  andx g0932(.a(n60), .b(n43), .O(n973));
  andx g0933(.a(n48), .b(n107), .O(n974));
  andx g0934(.a(n974), .b(n973), .O(n975));
  andx g0935(.a(n681), .b(n364), .O(n976));
  andx g0936(.a(n976), .b(n138), .O(n977));
  andx g0937(.a(n459), .b(n56), .O(n978));
  andx g0938(.a(n855), .b(n679), .O(n979));
  andx g0939(.a(n979), .b(n978), .O(n980));
  andx g0940(.a(n980), .b(n977), .O(n981));
  andx g0941(.a(n981), .b(n975), .O(n982));
  andx g0942(.a(n814), .b(n75), .O(n983));
  andx g0943(.a(n770), .b(n204), .O(n984));
  andx g0944(.a(n164), .b(n58), .O(n985));
  andx g0945(.a(n855), .b(n343), .O(n986));
  andx g0946(.a(n986), .b(n985), .O(n987));
  andx g0947(.a(n987), .b(n984), .O(n988));
  andx g0948(.a(n988), .b(n983), .O(n989));
  orx  g0949(.a(n989), .b(n982), .O(n990));
  orx  g0950(.a(n990), .b(n972), .O(n991));
  orx  g0951(.a(n991), .b(n965), .O(n992));
  orx  g0952(.a(n992), .b(n942), .O(n993));
  andx g0953(.a(n428), .b(n349), .O(n994));
  andx g0954(.a(n88), .b(pi27), .O(n995));
  andx g0955(.a(n995), .b(n994), .O(n996));
  andx g0956(.a(n80), .b(n99), .O(n997));
  andx g0957(.a(n997), .b(n53), .O(n998));
  andx g0958(.a(n998), .b(n996), .O(n999));
  andx g0959(.a(n168), .b(pi11), .O(n1000));
  andx g0960(.a(n566), .b(n66), .O(n1001));
  andx g0961(.a(n431), .b(n149), .O(n1002));
  andx g0962(.a(n1002), .b(n1001), .O(n1003));
  andx g0963(.a(n1003), .b(n1000), .O(n1004));
  orx  g0964(.a(n1004), .b(n999), .O(n1005));
  andx g0965(.a(n432), .b(n63), .O(n1006));
  andx g0966(.a(n618), .b(n250), .O(n1007));
  andx g0967(.a(n358), .b(n329), .O(n1008));
  andx g0968(.a(n1008), .b(n1007), .O(n1009));
  andx g0969(.a(n1009), .b(n1006), .O(n1010));
  andx g0970(.a(n1010), .b(n429), .O(n1011));
  andx g0971(.a(n943), .b(n731), .O(n1012));
  andx g0972(.a(n268), .b(n56), .O(n1013));
  andx g0973(.a(n318), .b(n61), .O(n1014));
  andx g0974(.a(n935), .b(n861), .O(n1015));
  andx g0975(.a(n1015), .b(n1014), .O(n1016));
  andx g0976(.a(n1016), .b(n1013), .O(n1017));
  andx g0977(.a(n1017), .b(n1012), .O(n1018));
  orx  g0978(.a(n1018), .b(n1011), .O(n1019));
  orx  g0979(.a(n1019), .b(n1005), .O(n1020));
  andx g0980(.a(n93), .b(n249), .O(n1021));
  andx g0981(.a(n1021), .b(n91), .O(n1022));
  andx g0982(.a(n1022), .b(n429), .O(n1023));
  andx g0983(.a(n304), .b(n64), .O(n1024));
  andx g0984(.a(n1024), .b(n433), .O(n1025));
  andx g0985(.a(n1025), .b(n1023), .O(n1026));
  andx g0986(.a(n902), .b(n690), .O(n1027));
  andx g0987(.a(n1027), .b(n179), .O(n1028));
  orx  g0988(.a(n1028), .b(n1026), .O(n1029));
  andx g0989(.a(pi07), .b(n99), .O(n1030));
  andx g0990(.a(n1030), .b(n432), .O(n1031));
  andx g0991(.a(n1031), .b(n996), .O(n1032));
  andx g0992(.a(n694), .b(n254), .O(n1033));
  andx g0993(.a(n1033), .b(n431), .O(n1034));
  andx g0994(.a(n1034), .b(n109), .O(n1035));
  orx  g0995(.a(n1035), .b(n1032), .O(n1036));
  orx  g0996(.a(n1036), .b(n1029), .O(n1037));
  orx  g0997(.a(n1037), .b(n1020), .O(n1038));
  andx g0998(.a(n484), .b(n91), .O(n1039));
  andx g0999(.a(n1039), .b(n145), .O(n1040));
  andx g1000(.a(n557), .b(n75), .O(n1041));
  andx g1001(.a(n1041), .b(n1040), .O(n1042));
  andx g1002(.a(n1042), .b(n818), .O(n1043));
  andx g1003(.a(n973), .b(n676), .O(n1044));
  andx g1004(.a(n120), .b(n68), .O(n1045));
  andx g1005(.a(n1045), .b(n897), .O(n1046));
  andx g1006(.a(n1046), .b(n1013), .O(n1047));
  andx g1007(.a(n1047), .b(n1044), .O(n1048));
  orx  g1008(.a(n1048), .b(n1043), .O(n1049));
  andx g1009(.a(n300), .b(n75), .O(n1050));
  andx g1010(.a(n536), .b(n323), .O(n1051));
  andx g1011(.a(n430), .b(n343), .O(n1052));
  andx g1012(.a(n1052), .b(n984), .O(n1053));
  andx g1013(.a(n1053), .b(n1051), .O(n1054));
  andx g1014(.a(n1054), .b(n1050), .O(n1055));
  andx g1015(.a(n973), .b(n48), .O(n1056));
  andx g1016(.a(n1056), .b(n42), .O(n1057));
  andx g1017(.a(n1057), .b(n301), .O(n1058));
  andx g1018(.a(n494), .b(n63), .O(n1059));
  andx g1019(.a(n307), .b(n254), .O(n1060));
  andx g1020(.a(n430), .b(n358), .O(n1061));
  andx g1021(.a(n1061), .b(n1060), .O(n1062));
  andx g1022(.a(n1062), .b(n1059), .O(n1063));
  andx g1023(.a(n1063), .b(n1058), .O(n1064));
  orx  g1024(.a(n1064), .b(n1055), .O(n1065));
  orx  g1025(.a(n1065), .b(n1049), .O(n1066));
  andx g1026(.a(n1027), .b(n83), .O(n1067));
  andx g1027(.a(n268), .b(n207), .O(n1068));
  andx g1028(.a(n1068), .b(n1014), .O(n1069));
  andx g1029(.a(n1069), .b(n1012), .O(n1070));
  orx  g1030(.a(n1070), .b(n1067), .O(n1071));
  andx g1031(.a(n566), .b(n50), .O(n1072));
  andx g1032(.a(n119), .b(n94), .O(n1073));
  andx g1033(.a(n536), .b(n343), .O(n1074));
  andx g1034(.a(n254), .b(n65), .O(n1075));
  andx g1035(.a(n1075), .b(n1074), .O(n1076));
  andx g1036(.a(n1076), .b(n1073), .O(n1077));
  andx g1037(.a(n1077), .b(n1072), .O(n1078));
  andx g1038(.a(pi34), .b(n99), .O(n1079));
  andx g1039(.a(pi29), .b(n87), .O(n1080));
  andx g1040(.a(n1080), .b(n229), .O(n1081));
  andx g1041(.a(n1081), .b(n1079), .O(n1082));
  andx g1042(.a(n1082), .b(n196), .O(n1083));
  orx  g1043(.a(n1083), .b(n1078), .O(n1084));
  orx  g1044(.a(n1084), .b(n1071), .O(n1085));
  orx  g1045(.a(n1085), .b(n1066), .O(n1086));
  orx  g1046(.a(n1086), .b(n1038), .O(n1087));
  orx  g1047(.a(n1087), .b(n993), .O(n1088));
  andx g1048(.a(n438), .b(n364), .O(n1089));
  andx g1049(.a(n756), .b(n119), .O(n1090));
  andx g1050(.a(n1090), .b(n1089), .O(n1091));
  andx g1051(.a(n1091), .b(n1051), .O(n1092));
  andx g1052(.a(n1092), .b(n1072), .O(n1093));
  andx g1053(.a(n213), .b(n214), .O(n1094));
  andx g1054(.a(n369), .b(n104), .O(n1095));
  andx g1055(.a(n494), .b(n304), .O(n1096));
  andx g1056(.a(n1096), .b(n1095), .O(n1097));
  andx g1057(.a(n1097), .b(n1094), .O(n1098));
  andx g1058(.a(n1098), .b(n732), .O(n1099));
  orx  g1059(.a(n1099), .b(n1093), .O(n1100));
  andx g1060(.a(n943), .b(n87), .O(n1101));
  andx g1061(.a(n127), .b(n101), .O(n1102));
  andx g1062(.a(n770), .b(n100), .O(n1103));
  andx g1063(.a(n679), .b(n204), .O(n1104));
  andx g1064(.a(n1104), .b(n1103), .O(n1105));
  andx g1065(.a(n1105), .b(n1102), .O(n1106));
  andx g1066(.a(n1106), .b(n1101), .O(n1107));
  andx g1067(.a(n494), .b(n364), .O(n1108));
  andx g1068(.a(n647), .b(n430), .O(n1109));
  andx g1069(.a(n307), .b(n101), .O(n1110));
  andx g1070(.a(n1110), .b(n1109), .O(n1111));
  andx g1071(.a(n1111), .b(n1108), .O(n1112));
  andx g1072(.a(n1112), .b(n983), .O(n1113));
  orx  g1073(.a(n1113), .b(n1107), .O(n1114));
  orx  g1074(.a(n1114), .b(n1100), .O(n1115));
  andx g1075(.a(n618), .b(n101), .O(n1116));
  andx g1076(.a(n1116), .b(n1042), .O(n1117));
  andx g1077(.a(n264), .b(n58), .O(n1118));
  andx g1078(.a(n818), .b(n1118), .O(n1119));
  andx g1079(.a(n1119), .b(n984), .O(n1120));
  andx g1080(.a(n1120), .b(n815), .O(n1121));
  orx  g1081(.a(n1121), .b(n1117), .O(n1122));
  andx g1082(.a(n756), .b(n66), .O(n1123));
  andx g1083(.a(n735), .b(n609), .O(n1124));
  andx g1084(.a(n1124), .b(n1123), .O(n1125));
  andx g1085(.a(n1125), .b(n169), .O(n1126));
  andx g1086(.a(n756), .b(n63), .O(n1127));
  andx g1087(.a(n1127), .b(n438), .O(n1128));
  andx g1088(.a(n1128), .b(n97), .O(n1129));
  orx  g1089(.a(n1129), .b(n1126), .O(n1130));
  orx  g1090(.a(n1130), .b(n1122), .O(n1131));
  orx  g1091(.a(n1131), .b(n1115), .O(n1132));
  andx g1092(.a(n369), .b(n171), .O(n1133));
  andx g1093(.a(n1133), .b(n682), .O(n1134));
  andx g1094(.a(n1134), .b(n807), .O(n1135));
  andx g1095(.a(n1135), .b(n1101), .O(n1136));
  andx g1096(.a(n818), .b(n264), .O(n1137));
  andx g1097(.a(n849), .b(n841), .O(n1138));
  andx g1098(.a(n1138), .b(n1137), .O(n1139));
  andx g1099(.a(n1139), .b(n814), .O(n1140));
  orx  g1100(.a(n1140), .b(n1136), .O(n1141));
  andx g1101(.a(n1057), .b(n88), .O(n1142));
  andx g1102(.a(n557), .b(n164), .O(n1143));
  andx g1103(.a(n304), .b(n254), .O(n1144));
  andx g1104(.a(n1144), .b(n1143), .O(n1145));
  andx g1105(.a(n1145), .b(n588), .O(n1146));
  andx g1106(.a(n1146), .b(n1142), .O(n1147));
  andx g1107(.a(n303), .b(n57), .O(n1148));
  andx g1108(.a(n1148), .b(n431), .O(n1149));
  andx g1109(.a(n661), .b(n1149), .O(n1150));
  andx g1110(.a(n1150), .b(n163), .O(n1151));
  andx g1111(.a(n1151), .b(n1058), .O(n1152));
  orx  g1112(.a(n1152), .b(n1147), .O(n1153));
  orx  g1113(.a(n1153), .b(n1141), .O(n1154));
  andx g1114(.a(n751), .b(n303), .O(n1155));
  andx g1115(.a(n944), .b(n250), .O(n1156));
  andx g1116(.a(n1156), .b(n1155), .O(n1157));
  andx g1117(.a(n1157), .b(n190), .O(n1158));
  andx g1118(.a(n860), .b(n829), .O(n1159));
  orx  g1119(.a(n1159), .b(n1158), .O(n1160));
  andx g1120(.a(n494), .b(n358), .O(n1161));
  andx g1121(.a(n1161), .b(n1095), .O(n1162));
  andx g1122(.a(n1162), .b(n1094), .O(n1163));
  andx g1123(.a(n1163), .b(n868), .O(n1164));
  andx g1124(.a(n90), .b(n212), .O(n1165));
  andx g1125(.a(n668), .b(n1165), .O(n1166));
  andx g1126(.a(n1166), .b(n639), .O(n1167));
  orx  g1127(.a(n1167), .b(n1164), .O(n1168));
  orx  g1128(.a(n1168), .b(n1160), .O(n1169));
  orx  g1129(.a(n1169), .b(n1154), .O(n1170));
  orx  g1130(.a(n1170), .b(n1132), .O(n1171));
  andx g1131(.a(n204), .b(n164), .O(n1172));
  andx g1132(.a(n1172), .b(n1144), .O(n1173));
  andx g1133(.a(n1173), .b(n894), .O(n1174));
  andx g1134(.a(n1174), .b(n893), .O(n1175));
  andx g1135(.a(n430), .b(n171), .O(n1176));
  andx g1136(.a(n1176), .b(n1110), .O(n1177));
  andx g1137(.a(n1177), .b(n577), .O(n1178));
  andx g1138(.a(n1178), .b(n302), .O(n1179));
  orx  g1139(.a(n1179), .b(n1175), .O(n1180));
  andx g1140(.a(n1109), .b(n418), .O(n1181));
  andx g1141(.a(n1181), .b(n1051), .O(n1182));
  andx g1142(.a(n1182), .b(n1050), .O(n1183));
  andx g1143(.a(n300), .b(n87), .O(n1184));
  andx g1144(.a(n984), .b(n489), .O(n1185));
  andx g1145(.a(n1185), .b(n1051), .O(n1186));
  andx g1146(.a(n1186), .b(n1184), .O(n1187));
  orx  g1147(.a(n1187), .b(n1183), .O(n1188));
  orx  g1148(.a(n1188), .b(n1180), .O(n1189));
  andx g1149(.a(n566), .b(pi29), .O(n1190));
  andx g1150(.a(n431), .b(n90), .O(n1191));
  andx g1151(.a(n1191), .b(n100), .O(n1192));
  andx g1152(.a(n1192), .b(n1190), .O(n1193));
  andx g1153(.a(n1193), .b(n717), .O(n1194));
  andx g1154(.a(n907), .b(n60), .O(n1195));
  andx g1155(.a(n909), .b(n431), .O(n1196));
  andx g1156(.a(n1196), .b(n100), .O(n1197));
  andx g1157(.a(n91), .b(n66), .O(n1198));
  andx g1158(.a(n1198), .b(n358), .O(n1199));
  andx g1159(.a(n1199), .b(n1197), .O(n1200));
  andx g1160(.a(n1200), .b(n1195), .O(n1201));
  orx  g1161(.a(n1201), .b(n1194), .O(n1202));
  andx g1162(.a(n781), .b(n751), .O(n1203));
  andx g1163(.a(n303), .b(n59), .O(n1204));
  andx g1164(.a(n1204), .b(n428), .O(n1205));
  andx g1165(.a(n1205), .b(n870), .O(n1206));
  andx g1166(.a(n1206), .b(n1203), .O(n1207));
  andx g1167(.a(n1207), .b(n975), .O(n1208));
  andx g1168(.a(n264), .b(n87), .O(n1209));
  andx g1169(.a(n1209), .b(n814), .O(n1210));
  andx g1170(.a(n935), .b(n214), .O(n1211));
  andx g1171(.a(n318), .b(n144), .O(n1212));
  andx g1172(.a(n430), .b(n104), .O(n1213));
  andx g1173(.a(n1213), .b(n1212), .O(n1214));
  andx g1174(.a(n1214), .b(n1211), .O(n1215));
  andx g1175(.a(n1215), .b(n1210), .O(n1216));
  orx  g1176(.a(n1216), .b(n1208), .O(n1217));
  orx  g1177(.a(n1217), .b(n1202), .O(n1218));
  orx  g1178(.a(n1218), .b(n1189), .O(n1219));
  andx g1179(.a(n536), .b(n144), .O(n1220));
  andx g1180(.a(n206), .b(n72), .O(n1221));
  andx g1181(.a(n1221), .b(n1220), .O(n1222));
  andx g1182(.a(n1222), .b(n968), .O(n1223));
  andx g1183(.a(n1223), .b(n300), .O(n1224));
  andx g1184(.a(n866), .b(n826), .O(n1225));
  orx  g1185(.a(n1225), .b(n1224), .O(n1226));
  andx g1186(.a(n90), .b(n57), .O(n1227));
  andx g1187(.a(n552), .b(n431), .O(n1228));
  andx g1188(.a(n618), .b(n264), .O(n1229));
  andx g1189(.a(n1229), .b(n1228), .O(n1230));
  andx g1190(.a(n1230), .b(n1227), .O(n1231));
  andx g1191(.a(n1231), .b(n1058), .O(n1232));
  andx g1192(.a(n171), .b(n101), .O(n1233));
  andx g1193(.a(n1233), .b(n1109), .O(n1234));
  andx g1194(.a(n1234), .b(n807), .O(n1235));
  andx g1195(.a(n1235), .b(n1184), .O(n1236));
  orx  g1196(.a(n1236), .b(n1232), .O(n1237));
  orx  g1197(.a(n1237), .b(n1226), .O(n1238));
  andx g1198(.a(n171), .b(n152), .O(n1239));
  andx g1199(.a(n1239), .b(n154), .O(n1240));
  andx g1200(.a(n1240), .b(n169), .O(n1241));
  andx g1201(.a(n48), .b(n56), .O(n1242));
  andx g1202(.a(n1242), .b(n45), .O(n1243));
  andx g1203(.a(n514), .b(n204), .O(n1244));
  andx g1204(.a(n264), .b(n120), .O(n1245));
  andx g1205(.a(n1245), .b(n1244), .O(n1246));
  andx g1206(.a(n1246), .b(n349), .O(n1247));
  andx g1207(.a(n1247), .b(n1243), .O(n1248));
  orx  g1208(.a(n1248), .b(n1241), .O(n1249));
  andx g1209(.a(n751), .b(n101), .O(n1250));
  andx g1210(.a(n1250), .b(n966), .O(n1251));
  andx g1211(.a(n117), .b(n101), .O(n1252));
  andx g1212(.a(n1252), .b(n870), .O(n1253));
  andx g1213(.a(n1253), .b(n470), .O(n1254));
  andx g1214(.a(n1254), .b(n1012), .O(n1255));
  orx  g1215(.a(n1255), .b(n1251), .O(n1256));
  orx  g1216(.a(n1256), .b(n1249), .O(n1257));
  orx  g1217(.a(n1257), .b(n1238), .O(n1258));
  orx  g1218(.a(n1258), .b(n1219), .O(n1259));
  orx  g1219(.a(n1259), .b(n1171), .O(n1260));
  orx  g1220(.a(n1260), .b(n1088), .O(n1261));
  andx g1221(.a(n369), .b(n337), .O(n1262));
  andx g1222(.a(n1262), .b(n336), .O(n1263));
  andx g1223(.a(n1263), .b(n335), .O(n1264));
  andx g1224(.a(pi17), .b(n212), .O(n1265));
  andx g1225(.a(n1265), .b(n104), .O(n1266));
  andx g1226(.a(n459), .b(n110), .O(n1267));
  andx g1227(.a(n1267), .b(n1266), .O(n1268));
  andx g1228(.a(n1268), .b(n638), .O(n1269));
  orx  g1229(.a(n1269), .b(n1264), .O(n1270));
  andx g1230(.a(pi34), .b(pi29), .O(n1271));
  andx g1231(.a(n1271), .b(n120), .O(n1272));
  andx g1232(.a(n1272), .b(n100), .O(n1273));
  andx g1233(.a(n1273), .b(n190), .O(n1274));
  andx g1234(.a(n438), .b(n397), .O(n1275));
  andx g1235(.a(n1275), .b(n1123), .O(n1276));
  andx g1236(.a(n1276), .b(n396), .O(n1277));
  orx  g1237(.a(n1277), .b(n1274), .O(n1278));
  orx  g1238(.a(n1278), .b(n1270), .O(n1279));
  andx g1239(.a(pi24), .b(n66), .O(n1280));
  andx g1240(.a(n431), .b(pi23), .O(n1281));
  andx g1241(.a(n1281), .b(n1280), .O(n1282));
  andx g1242(.a(n1282), .b(n256), .O(n1283));
  andx g1243(.a(n62), .b(n92), .O(n1284));
  andx g1244(.a(n960), .b(n690), .O(n1285));
  andx g1245(.a(n1285), .b(n1284), .O(n1286));
  orx  g1246(.a(n1286), .b(n1283), .O(n1287));
  andx g1247(.a(n749), .b(n198), .O(n1288));
  andx g1248(.a(n1288), .b(n274), .O(n1289));
  andx g1249(.a(n292), .b(n108), .O(n1290));
  andx g1250(.a(n1290), .b(n1289), .O(n1291));
  andx g1251(.a(n1198), .b(n264), .O(n1292));
  andx g1252(.a(n42), .b(n249), .O(n1293));
  andx g1253(.a(n1293), .b(n267), .O(n1294));
  andx g1254(.a(n1294), .b(n1292), .O(n1295));
  andx g1255(.a(n304), .b(n63), .O(n1296));
  andx g1256(.a(n1296), .b(n62), .O(n1297));
  andx g1257(.a(n1297), .b(n1295), .O(n1298));
  orx  g1258(.a(n1298), .b(n1291), .O(n1299));
  orx  g1259(.a(n1299), .b(n1287), .O(n1300));
  orx  g1260(.a(n1300), .b(n1279), .O(n1301));
  andx g1261(.a(n358), .b(n345), .O(n1302));
  andx g1262(.a(n1302), .b(n200), .O(n1303));
  andx g1263(.a(n1303), .b(n342), .O(n1304));
  andx g1264(.a(n431), .b(n66), .O(n1305));
  andx g1265(.a(n1305), .b(n661), .O(n1306));
  andx g1266(.a(n1306), .b(n1284), .O(n1307));
  orx  g1267(.a(n1307), .b(n1304), .O(n1308));
  andx g1268(.a(n287), .b(n234), .O(n1309));
  andx g1269(.a(n238), .b(n58), .O(n1310));
  andx g1270(.a(n1310), .b(n241), .O(n1311));
  andx g1271(.a(n1311), .b(n237), .O(n1312));
  orx  g1272(.a(n1312), .b(n1309), .O(n1313));
  orx  g1273(.a(n1313), .b(n1308), .O(n1314));
  andx g1274(.a(pi25), .b(n60), .O(n1315));
  andx g1275(.a(n1315), .b(n88), .O(n1316));
  andx g1276(.a(n1316), .b(n117), .O(n1317));
  andx g1277(.a(n1280), .b(n199), .O(n1318));
  andx g1278(.a(n1318), .b(n756), .O(n1319));
  andx g1279(.a(n1319), .b(n1317), .O(n1320));
  andx g1280(.a(n313), .b(n144), .O(n1321));
  andx g1281(.a(n91), .b(n57), .O(n1322));
  andx g1282(.a(n1322), .b(n318), .O(n1323));
  andx g1283(.a(n1323), .b(n1321), .O(n1324));
  andx g1284(.a(n1324), .b(n1197), .O(n1325));
  orx  g1285(.a(n1325), .b(n1320), .O(n1326));
  andx g1286(.a(n120), .b(n81), .O(n1327));
  andx g1287(.a(n1327), .b(n1006), .O(n1328));
  andx g1288(.a(n1328), .b(n792), .O(n1329));
  andx g1289(.a(n1198), .b(n138), .O(n1330));
  andx g1290(.a(n909), .b(n267), .O(n1331));
  andx g1291(.a(n1331), .b(n1330), .O(n1332));
  andx g1292(.a(n60), .b(n93), .O(n1333));
  andx g1293(.a(n1333), .b(n58), .O(n1334));
  andx g1294(.a(n855), .b(n249), .O(n1335));
  andx g1295(.a(n1335), .b(n1334), .O(n1336));
  andx g1296(.a(n1336), .b(n1332), .O(n1337));
  orx  g1297(.a(n1337), .b(n1329), .O(n1338));
  orx  g1298(.a(n1338), .b(n1326), .O(n1339));
  orx  g1299(.a(n1339), .b(n1314), .O(n1340));
  orx  g1300(.a(n1340), .b(n1301), .O(n1341));
  andx g1301(.a(n429), .b(n92), .O(n1342));
  andx g1302(.a(n164), .b(n63), .O(n1343));
  andx g1303(.a(n75), .b(n87), .O(n1344));
  andx g1304(.a(n1344), .b(n523), .O(n1345));
  andx g1305(.a(n1345), .b(n1343), .O(n1346));
  andx g1306(.a(n1346), .b(n1342), .O(n1347));
  andx g1307(.a(n922), .b(n94), .O(n1348));
  andx g1308(.a(n855), .b(n718), .O(n1349));
  andx g1309(.a(n99), .b(n249), .O(n1350));
  andx g1310(.a(n1350), .b(n204), .O(n1351));
  andx g1311(.a(n1351), .b(n944), .O(n1352));
  andx g1312(.a(n1352), .b(n1349), .O(n1353));
  andx g1313(.a(n1353), .b(n1348), .O(n1354));
  orx  g1314(.a(n1354), .b(n1347), .O(n1355));
  andx g1315(.a(n892), .b(n88), .O(n1356));
  andx g1316(.a(n249), .b(n66), .O(n1357));
  andx g1317(.a(n1357), .b(n895), .O(n1358));
  andx g1318(.a(n1345), .b(n1358), .O(n1359));
  andx g1319(.a(n1359), .b(n712), .O(n1360));
  andx g1320(.a(n1360), .b(n1356), .O(n1361));
  andx g1321(.a(n1334), .b(n44), .O(n1362));
  andx g1322(.a(n1362), .b(n91), .O(n1363));
  andx g1323(.a(n318), .b(n53), .O(n1364));
  andx g1324(.a(n1364), .b(n712), .O(n1365));
  andx g1325(.a(n1365), .b(n1363), .O(n1366));
  orx  g1326(.a(n1366), .b(n1361), .O(n1367));
  orx  g1327(.a(n1367), .b(n1355), .O(n1368));
  andx g1328(.a(n557), .b(n358), .O(n1369));
  andx g1329(.a(n855), .b(n269), .O(n1370));
  andx g1330(.a(n1370), .b(n449), .O(n1371));
  andx g1331(.a(n1371), .b(n1369), .O(n1372));
  andx g1332(.a(n376), .b(n231), .O(n1373));
  orx  g1333(.a(n1373), .b(n1372), .O(n1374));
  andx g1334(.a(n861), .b(n404), .O(n1375));
  andx g1335(.a(n1375), .b(n144), .O(n1376));
  andx g1336(.a(n99), .b(n212), .O(n1377));
  andx g1337(.a(n1377), .b(n274), .O(n1378));
  andx g1338(.a(n1378), .b(n864), .O(n1379));
  andx g1339(.a(n1379), .b(n1376), .O(n1380));
  andx g1340(.a(n437), .b(pi28), .O(n1381));
  andx g1341(.a(n1381), .b(n264), .O(n1382));
  andx g1342(.a(n250), .b(n87), .O(n1383));
  andx g1343(.a(n1383), .b(n248), .O(n1384));
  andx g1344(.a(n1384), .b(n1382), .O(n1385));
  orx  g1345(.a(n1385), .b(n1380), .O(n1386));
  orx  g1346(.a(n1386), .b(n1374), .O(n1387));
  andx g1347(.a(pi30), .b(n67), .O(n1388));
  andx g1348(.a(n269), .b(n249), .O(n1389));
  andx g1349(.a(n1389), .b(n1388), .O(n1390));
  andx g1350(.a(n1390), .b(n1081), .O(n1391));
  andx g1351(.a(pi07), .b(pi27), .O(n1392));
  andx g1352(.a(n1392), .b(n250), .O(n1393));
  andx g1353(.a(n945), .b(n268), .O(n1394));
  andx g1354(.a(n1394), .b(n264), .O(n1395));
  andx g1355(.a(n1395), .b(n1393), .O(n1396));
  orx  g1356(.a(n1396), .b(n1391), .O(n1397));
  andx g1357(.a(pi25), .b(n67), .O(n1398));
  andx g1358(.a(n257), .b(n250), .O(n1399));
  andx g1359(.a(n1399), .b(n1398), .O(n1400));
  andx g1360(.a(n1400), .b(n1075), .O(n1401));
  andx g1361(.a(n388), .b(n234), .O(n1402));
  orx  g1362(.a(n1402), .b(n1401), .O(n1403));
  orx  g1363(.a(n1403), .b(n1397), .O(n1404));
  orx  g1364(.a(n1404), .b(n1387), .O(n1405));
  orx  g1365(.a(n1405), .b(n1368), .O(n1406));
  orx  g1366(.a(n1406), .b(n1341), .O(n1407));
  andx g1367(.a(n566), .b(n229), .O(n1408));
  andx g1368(.a(n1408), .b(n1327), .O(n1409));
  andx g1369(.a(n1409), .b(n146), .O(n1410));
  andx g1370(.a(n75), .b(pi24), .O(n1411));
  andx g1371(.a(n1411), .b(n250), .O(n1412));
  andx g1372(.a(n756), .b(n431), .O(n1413));
  andx g1373(.a(n1413), .b(n1398), .O(n1414));
  andx g1374(.a(n1414), .b(n1412), .O(n1415));
  orx  g1375(.a(n1415), .b(n1410), .O(n1416));
  andx g1376(.a(n449), .b(n257), .O(n1417));
  andx g1377(.a(n1417), .b(n72), .O(n1418));
  andx g1378(.a(n1418), .b(n1317), .O(n1419));
  andx g1379(.a(n660), .b(n66), .O(n1420));
  andx g1380(.a(n433), .b(n1420), .O(n1421));
  andx g1381(.a(n1421), .b(n396), .O(n1422));
  orx  g1382(.a(n1422), .b(n1419), .O(n1423));
  orx  g1383(.a(n1423), .b(n1416), .O(n1424));
  andx g1384(.a(n397), .b(n110), .O(n1425));
  andx g1385(.a(n1425), .b(n120), .O(n1426));
  andx g1386(.a(n1426), .b(n665), .O(n1427));
  andx g1387(.a(n120), .b(n72), .O(n1428));
  andx g1388(.a(n1428), .b(n110), .O(n1429));
  andx g1389(.a(n1429), .b(n178), .O(n1430));
  orx  g1390(.a(n1430), .b(n1427), .O(n1431));
  andx g1391(.a(n1315), .b(n56), .O(n1432));
  andx g1392(.a(n1432), .b(n76), .O(n1433));
  andx g1393(.a(n1433), .b(n1418), .O(n1434));
  andx g1394(.a(n388), .b(n284), .O(n1435));
  orx  g1395(.a(n1435), .b(n1434), .O(n1436));
  orx  g1396(.a(n1436), .b(n1431), .O(n1437));
  orx  g1397(.a(n1437), .b(n1424), .O(n1438));
  andx g1398(.a(n902), .b(n52), .O(n1439));
  andx g1399(.a(n1439), .b(n358), .O(n1440));
  andx g1400(.a(n1440), .b(n658), .O(n1441));
  andx g1401(.a(pi24), .b(n249), .O(n1442));
  andx g1402(.a(pi23), .b(n67), .O(n1443));
  andx g1403(.a(n1443), .b(n1442), .O(n1444));
  andx g1404(.a(n1344), .b(n269), .O(n1445));
  andx g1405(.a(n1445), .b(n65), .O(n1446));
  andx g1406(.a(n1446), .b(n1444), .O(n1447));
  orx  g1407(.a(n1447), .b(n1441), .O(n1448));
  andx g1408(.a(n204), .b(n117), .O(n1449));
  andx g1409(.a(n1449), .b(n855), .O(n1450));
  andx g1410(.a(n250), .b(n120), .O(n1451));
  andx g1411(.a(n1451), .b(n752), .O(n1452));
  andx g1412(.a(n1452), .b(n1450), .O(n1453));
  andx g1413(.a(n75), .b(n91), .O(n1454));
  andx g1414(.a(n1454), .b(pi25), .O(n1455));
  andx g1415(.a(n1455), .b(n1442), .O(n1456));
  andx g1416(.a(n1456), .b(n247), .O(n1457));
  orx  g1417(.a(n1457), .b(n1453), .O(n1458));
  orx  g1418(.a(n1458), .b(n1448), .O(n1459));
  andx g1419(.a(n1080), .b(n1079), .O(n1460));
  andx g1420(.a(n1460), .b(n432), .O(n1461));
  andx g1421(.a(n1461), .b(n700), .O(n1462));
  andx g1422(.a(n855), .b(n250), .O(n1463));
  andx g1423(.a(n432), .b(n329), .O(n1464));
  andx g1424(.a(n1464), .b(n1463), .O(n1465));
  andx g1425(.a(n514), .b(n66), .O(n1466));
  andx g1426(.a(n1466), .b(n137), .O(n1467));
  andx g1427(.a(n1467), .b(n1465), .O(n1468));
  orx  g1428(.a(n1468), .b(n1462), .O(n1469));
  andx g1429(.a(n358), .b(n73), .O(n1470));
  andx g1430(.a(n1470), .b(n286), .O(n1471));
  andx g1431(.a(n1471), .b(n1284), .O(n1472));
  andx g1432(.a(n200), .b(n245), .O(n1473));
  andx g1433(.a(n250), .b(n248), .O(n1474));
  andx g1434(.a(n1474), .b(n1473), .O(n1475));
  orx  g1435(.a(n1475), .b(n1472), .O(n1476));
  orx  g1436(.a(n1476), .b(n1469), .O(n1477));
  orx  g1437(.a(n1477), .b(n1459), .O(n1478));
  orx  g1438(.a(n1478), .b(n1438), .O(n1479));
  andx g1439(.a(n450), .b(n110), .O(n1480));
  andx g1440(.a(n1480), .b(n129), .O(n1481));
  andx g1441(.a(n292), .b(n1327), .O(n1482));
  andx g1442(.a(n1482), .b(n217), .O(n1483));
  orx  g1443(.a(n1483), .b(n1481), .O(n1484));
  andx g1444(.a(pi36), .b(n249), .O(n1485));
  andx g1445(.a(n1485), .b(n264), .O(n1486));
  andx g1446(.a(n603), .b(n92), .O(n1487));
  andx g1447(.a(n1487), .b(n1486), .O(n1488));
  andx g1448(.a(n386), .b(n231), .O(n1489));
  orx  g1449(.a(n1489), .b(n1488), .O(n1490));
  orx  g1450(.a(n1490), .b(n1484), .O(n1491));
  andx g1451(.a(n149), .b(n130), .O(n1492));
  andx g1452(.a(n1492), .b(n1305), .O(n1493));
  andx g1453(.a(n1493), .b(n79), .O(n1494));
  andx g1454(.a(n304), .b(n250), .O(n1495));
  andx g1455(.a(n182), .b(n104), .O(n1496));
  andx g1456(.a(n1496), .b(n164), .O(n1497));
  andx g1457(.a(n1497), .b(n1495), .O(n1498));
  orx  g1458(.a(n1498), .b(n1494), .O(n1499));
  andx g1459(.a(n1079), .b(n432), .O(n1500));
  andx g1460(.a(n1500), .b(n120), .O(n1501));
  andx g1461(.a(n1501), .b(n994), .O(n1502));
  andx g1462(.a(n91), .b(n87), .O(n1503));
  andx g1463(.a(n1503), .b(pi25), .O(n1504));
  andx g1464(.a(n1504), .b(n1442), .O(n1505));
  andx g1465(.a(n1505), .b(n1382), .O(n1506));
  orx  g1466(.a(n1506), .b(n1502), .O(n1507));
  orx  g1467(.a(n1507), .b(n1499), .O(n1508));
  orx  g1468(.a(n1508), .b(n1491), .O(n1509));
  andx g1469(.a(n545), .b(n63), .O(n1510));
  andx g1470(.a(n357), .b(n138), .O(n1511));
  andx g1471(.a(n1511), .b(n1510), .O(n1512));
  andx g1472(.a(n1512), .b(n1040), .O(n1513));
  andx g1473(.a(n53), .b(pi24), .O(n1514));
  andx g1474(.a(n1514), .b(n1443), .O(n1515));
  andx g1475(.a(n1515), .b(n379), .O(n1516));
  orx  g1476(.a(n1516), .b(n1513), .O(n1517));
  andx g1477(.a(n334), .b(n254), .O(n1518));
  andx g1478(.a(n273), .b(n72), .O(n1519));
  andx g1479(.a(n1519), .b(n1518), .O(n1520));
  andx g1480(.a(n1520), .b(n403), .O(n1521));
  andx g1481(.a(n388), .b(n386), .O(n1522));
  orx  g1482(.a(n1522), .b(n1521), .O(n1523));
  orx  g1483(.a(n1523), .b(n1517), .O(n1524));
  andx g1484(.a(n164), .b(pi07), .O(n1525));
  andx g1485(.a(n1525), .b(n138), .O(n1526));
  andx g1486(.a(n1526), .b(n658), .O(n1527));
  andx g1487(.a(pi30), .b(pi29), .O(n1528));
  andx g1488(.a(n381), .b(n52), .O(n1529));
  andx g1489(.a(n1529), .b(n1528), .O(n1530));
  andx g1490(.a(n1530), .b(n378), .O(n1531));
  orx  g1491(.a(n1531), .b(n1527), .O(n1532));
  andx g1492(.a(n1319), .b(n1433), .O(n1533));
  andx g1493(.a(pi25), .b(pi24), .O(n1534));
  andx g1494(.a(n1534), .b(n250), .O(n1535));
  andx g1495(.a(n1535), .b(n1473), .O(n1536));
  orx  g1496(.a(n1536), .b(n1533), .O(n1537));
  orx  g1497(.a(n1537), .b(n1532), .O(n1538));
  orx  g1498(.a(n1538), .b(n1524), .O(n1539));
  orx  g1499(.a(n1539), .b(n1509), .O(n1540));
  orx  g1500(.a(n1540), .b(n1479), .O(n1541));
  orx  g1501(.a(n1541), .b(n1407), .O(n1542));
  andx g1502(.a(n878), .b(n667), .O(n1543));
  andx g1503(.a(n254), .b(n56), .O(n1544));
  andx g1504(.a(n2665), .b(n80), .O(n1545));
  andx g1505(.a(n1545), .b(n1282), .O(n1546));
  orx  g1506(.a(n1546), .b(n1543), .O(n1547));
  andx g1507(.a(n182), .b(n65), .O(n1548));
  andx g1508(.a(n1548), .b(n667), .O(n1549));
  andx g1509(.a(n343), .b(n171), .O(n1550));
  andx g1510(.a(n1550), .b(n712), .O(n1551));
  andx g1511(.a(n1551), .b(n1363), .O(n1552));
  orx  g1512(.a(n1552), .b(n1549), .O(n1553));
  orx  g1513(.a(n1553), .b(n1547), .O(n1554));
  andx g1514(.a(n609), .b(n63), .O(n1555));
  andx g1515(.a(n784), .b(n152), .O(n1556));
  andx g1516(.a(n1556), .b(n1555), .O(n1557));
  andx g1517(.a(n1557), .b(n148), .O(n1558));
  andx g1518(.a(n878), .b(n795), .O(n1559));
  orx  g1519(.a(n1559), .b(n1558), .O(n1560));
  andx g1520(.a(n459), .b(n138), .O(n1561));
  andx g1521(.a(n1561), .b(n712), .O(n1562));
  andx g1522(.a(n1562), .b(n1363), .O(n1563));
  andx g1523(.a(n1333), .b(n922), .O(n1564));
  andx g1524(.a(n1564), .b(n88), .O(n1565));
  andx g1525(.a(n1485), .b(n718), .O(n1566));
  andx g1526(.a(n1344), .b(n618), .O(n1567));
  andx g1527(.a(n1567), .b(n1566), .O(n1568));
  andx g1528(.a(n1568), .b(n588), .O(n1569));
  andx g1529(.a(n1569), .b(n1565), .O(n1570));
  orx  g1530(.a(n1570), .b(n1563), .O(n1571));
  orx  g1531(.a(n1571), .b(n1560), .O(n1572));
  orx  g1532(.a(n1572), .b(n1554), .O(n1573));
  andx g1533(.a(n1545), .b(n260), .O(n1574));
  andx g1534(.a(n995), .b(n190), .O(n1575));
  andx g1535(.a(n1575), .b(n710), .O(n1576));
  orx  g1536(.a(n1576), .b(n1574), .O(n1577));
  andx g1537(.a(n766), .b(n398), .O(n1578));
  andx g1538(.a(n1578), .b(n1023), .O(n1579));
  andx g1539(.a(n208), .b(n238), .O(n1580));
  andx g1540(.a(n1580), .b(n629), .O(n1581));
  andx g1541(.a(n1581), .b(n468), .O(n1582));
  orx  g1542(.a(n1582), .b(n1579), .O(n1583));
  orx  g1543(.a(n1583), .b(n1577), .O(n1584));
  andx g1544(.a(n193), .b(n120), .O(n1585));
  andx g1545(.a(n1585), .b(n191), .O(n1586));
  andx g1546(.a(n691), .b(n131), .O(n1587));
  orx  g1547(.a(n1587), .b(n1586), .O(n1588));
  andx g1548(.a(n1575), .b(n706), .O(n1589));
  andx g1549(.a(n1027), .b(n131), .O(n1590));
  orx  g1550(.a(n1590), .b(n1589), .O(n1591));
  orx  g1551(.a(n1591), .b(n1588), .O(n1592));
  orx  g1552(.a(n1592), .b(n1584), .O(n1593));
  orx  g1553(.a(n1593), .b(n1573), .O(n1594));
  andx g1554(.a(n681), .b(n138), .O(n1595));
  andx g1555(.a(n1595), .b(n856), .O(n1596));
  andx g1556(.a(n1596), .b(n680), .O(n1597));
  andx g1557(.a(n1597), .b(n769), .O(n1598));
  andx g1558(.a(n1204), .b(n357), .O(n1599));
  andx g1559(.a(n1599), .b(n852), .O(n1600));
  andx g1560(.a(n1600), .b(n588), .O(n1601));
  andx g1561(.a(n1601), .b(n1142), .O(n1602));
  orx  g1562(.a(n1602), .b(n1598), .O(n1603));
  andx g1563(.a(n104), .b(n57), .O(n1604));
  andx g1564(.a(n264), .b(n204), .O(n1605));
  andx g1565(.a(n1605), .b(n1052), .O(n1606));
  andx g1566(.a(n1606), .b(n1604), .O(n1607));
  andx g1567(.a(n1607), .b(n893), .O(n1608));
  andx g1568(.a(n922), .b(n117), .O(n1609));
  andx g1569(.a(n303), .b(n66), .O(n1610));
  andx g1570(.a(n1610), .b(n198), .O(n1611));
  andx g1571(.a(n397), .b(n120), .O(n1612));
  andx g1572(.a(n1612), .b(n1486), .O(n1613));
  andx g1573(.a(n1613), .b(n1611), .O(n1614));
  andx g1574(.a(n1614), .b(n1609), .O(n1615));
  orx  g1575(.a(n1615), .b(n1608), .O(n1616));
  orx  g1576(.a(n1616), .b(n1603), .O(n1617));
  andx g1577(.a(n323), .b(n60), .O(n1618));
  andx g1578(.a(n1357), .b(n206), .O(n1619));
  andx g1579(.a(n1619), .b(n489), .O(n1620));
  andx g1580(.a(n1620), .b(n1618), .O(n1621));
  andx g1581(.a(n1621), .b(n543), .O(n1622));
  andx g1582(.a(n1233), .b(n545), .O(n1623));
  andx g1583(.a(n1623), .b(n937), .O(n1624));
  andx g1584(.a(n1624), .b(n300), .O(n1625));
  orx  g1585(.a(n1625), .b(n1622), .O(n1626));
  andx g1586(.a(pi26), .b(n107), .O(n1627));
  andx g1587(.a(n1627), .b(n922), .O(n1628));
  andx g1588(.a(n751), .b(n523), .O(n1629));
  andx g1589(.a(n1629), .b(n1344), .O(n1630));
  andx g1590(.a(n979), .b(n163), .O(n1631));
  andx g1591(.a(n1631), .b(n1630), .O(n1632));
  andx g1592(.a(n1632), .b(n1628), .O(n1633));
  andx g1593(.a(pi26), .b(n93), .O(n1634));
  andx g1594(.a(n1634), .b(n428), .O(n1635));
  andx g1595(.a(n902), .b(n536), .O(n1636));
  andx g1596(.a(n238), .b(n104), .O(n1637));
  andx g1597(.a(n1637), .b(n1636), .O(n1638));
  andx g1598(.a(n1638), .b(n1635), .O(n1639));
  andx g1599(.a(n1639), .b(n115), .O(n1640));
  orx  g1600(.a(n1640), .b(n1633), .O(n1641));
  orx  g1601(.a(n1641), .b(n1626), .O(n1642));
  orx  g1602(.a(n1642), .b(n1617), .O(n1643));
  andx g1603(.a(n795), .b(n670), .O(n1644));
  andx g1604(.a(n1357), .b(n343), .O(n1645));
  andx g1605(.a(n895), .b(n432), .O(n1646));
  andx g1606(.a(n1646), .b(n1645), .O(n1647));
  andx g1607(.a(n1647), .b(n712), .O(n1648));
  andx g1608(.a(n1648), .b(n1356), .O(n1649));
  orx  g1609(.a(n1649), .b(n1644), .O(n1650));
  andx g1610(.a(n922), .b(n144), .O(n1651));
  andx g1611(.a(n1651), .b(n88), .O(n1652));
  andx g1612(.a(n1344), .b(n514), .O(n1653));
  andx g1613(.a(n1653), .b(n1358), .O(n1654));
  andx g1614(.a(n1654), .b(n349), .O(n1655));
  andx g1615(.a(n1655), .b(n1652), .O(n1656));
  andx g1616(.a(n358), .b(n238), .O(n1657));
  andx g1617(.a(n1657), .b(n903), .O(n1658));
  andx g1618(.a(n1658), .b(n1342), .O(n1659));
  orx  g1619(.a(n1659), .b(n1656), .O(n1660));
  orx  g1620(.a(n1660), .b(n1650), .O(n1661));
  andx g1621(.a(n1204), .b(n491), .O(n1662));
  andx g1622(.a(n1662), .b(n1511), .O(n1663));
  andx g1623(.a(n1663), .b(n588), .O(n1664));
  andx g1624(.a(n1664), .b(n543), .O(n1665));
  andx g1625(.a(n494), .b(n60), .O(n1666));
  andx g1626(.a(n589), .b(n566), .O(n1667));
  andx g1627(.a(n1667), .b(n928), .O(n1668));
  andx g1628(.a(n1668), .b(n1666), .O(n1669));
  andx g1629(.a(n1669), .b(n1210), .O(n1670));
  orx  g1630(.a(n1670), .b(n1665), .O(n1671));
  andx g1631(.a(n523), .b(n264), .O(n1672));
  andx g1632(.a(n1672), .b(n522), .O(n1673));
  andx g1633(.a(n1673), .b(n1342), .O(n1674));
  andx g1634(.a(n1548), .b(n795), .O(n1675));
  orx  g1635(.a(n1675), .b(n1674), .O(n1676));
  orx  g1636(.a(n1676), .b(n1671), .O(n1677));
  orx  g1637(.a(n1677), .b(n1661), .O(n1678));
  orx  g1638(.a(n1678), .b(n1643), .O(n1679));
  orx  g1639(.a(n1679), .b(n1594), .O(n1680));
  orx  g1640(.a(n1680), .b(n1542), .O(n1681));
  orx  g1641(.a(n1681), .b(n1261), .O(n1682));
  orx  g1642(.a(n1682), .b(n884), .O(n1683));
  orx  g1643(.a(n1683), .b(n637), .O(po0));
  andx g1644(.a(n545), .b(pi37), .O(n1685));
  andx g1645(.a(n1454), .b(n104), .O(n1686));
  invx g1646(.a(pi24), .O(n1687));
  andx g1647(.a(n1687), .b(n64), .O(n1688));
  andx g1648(.a(n67), .b(n249), .O(n1689));
  andx g1649(.a(n1689), .b(n1688), .O(n1690));
  andx g1650(.a(n1690), .b(n1686), .O(n1691));
  andx g1651(.a(n1691), .b(n1685), .O(n1692));
  orx  g1652(.a(n1692), .b(n362), .O(n1693));
  andx g1653(.a(pi37), .b(n59), .O(n1694));
  invx g1654(.a(pi34), .O(n1695));
  andx g1655(.a(n1695), .b(n1687), .O(n1696));
  andx g1656(.a(n1696), .b(n1694), .O(n1697));
  andx g1657(.a(n1198), .b(n855), .O(n1698));
  andx g1658(.a(n1698), .b(n1697), .O(n1699));
  andx g1659(.a(n1344), .b(n277), .O(n1700));
  andx g1660(.a(n1700), .b(n1334), .O(n1701));
  andx g1661(.a(n1701), .b(n1699), .O(n1702));
  orx  g1662(.a(n1702), .b(n1435), .O(n1703));
  orx  g1663(.a(n1703), .b(n1693), .O(n1704));
  andx g1664(.a(n699), .b(n171), .O(n1705));
  andx g1665(.a(pi07), .b(n63), .O(n1706));
  andx g1666(.a(n595), .b(n289), .O(n1707));
  andx g1667(.a(n1707), .b(n1705), .O(n1708));
  orx  g1668(.a(n1708), .b(n387), .O(n1709));
  andx g1669(.a(n333), .b(pi28), .O(n1710));
  andx g1670(.a(n1710), .b(n58), .O(n1711));
  andx g1671(.a(n459), .b(n59), .O(n1712));
  andx g1672(.a(n404), .b(n397), .O(n1713));
  andx g1673(.a(n1713), .b(n1712), .O(n1714));
  andx g1674(.a(n1714), .b(n1711), .O(n1715));
  orx  g1675(.a(n1715), .b(n282), .O(n1716));
  orx  g1676(.a(n1716), .b(n1709), .O(n1717));
  orx  g1677(.a(n1717), .b(n1704), .O(n1718));
  andx g1678(.a(n250), .b(pi07), .O(n1719));
  andx g1679(.a(n67), .b(pi29), .O(n1720));
  andx g1680(.a(n254), .b(n220), .O(n1721));
  andx g1681(.a(n1721), .b(n1720), .O(n1722));
  andx g1682(.a(n1722), .b(n1719), .O(n1723));
  andx g1683(.a(n199), .b(n80), .O(n1724));
  andx g1684(.a(pi10), .b(pi11), .O(n1725));
  andx g1685(.a(n1725), .b(n756), .O(n1726));
  andx g1686(.a(n1726), .b(n1724), .O(n1727));
  andx g1687(.a(n1727), .b(n429), .O(n1728));
  orx  g1688(.a(n1728), .b(n1723), .O(n1729));
  andx g1689(.a(pi27), .b(n91), .O(n1730));
  andx g1690(.a(n1730), .b(n1689), .O(n1731));
  andx g1691(.a(pi24), .b(n63), .O(n1732));
  andx g1692(.a(pi23), .b(n52), .O(n1733));
  andx g1693(.a(n1733), .b(n1344), .O(n1734));
  andx g1694(.a(n1734), .b(n1732), .O(n1735));
  andx g1695(.a(n1735), .b(n1731), .O(n1736));
  orx  g1696(.a(n1736), .b(n1489), .O(n1737));
  orx  g1697(.a(n1737), .b(n1729), .O(n1738));
  orx  g1698(.a(n389), .b(n377), .O(n1739));
  andx g1699(.a(n88), .b(pi29), .O(n1740));
  andx g1700(.a(n1740), .b(n52), .O(n1741));
  andx g1701(.a(n1741), .b(n584), .O(n1742));
  andx g1702(.a(n1742), .b(n190), .O(n1743));
  orx  g1703(.a(n1743), .b(n1447), .O(n1744));
  orx  g1704(.a(n1744), .b(n1739), .O(n1745));
  orx  g1705(.a(n1745), .b(n1738), .O(n1746));
  orx  g1706(.a(n1746), .b(n1718), .O(n1747));
  andx g1707(.a(n53), .b(pi29), .O(n1748));
  andx g1708(.a(n1748), .b(n289), .O(n1749));
  andx g1709(.a(n1749), .b(n700), .O(n1750));
  andx g1710(.a(n254), .b(n144), .O(n1751));
  andx g1711(.a(n1751), .b(n1725), .O(n1752));
  andx g1712(.a(n88), .b(n66), .O(n1753));
  andx g1713(.a(n1428), .b(n1752), .O(n1754));
  orx  g1714(.a(n1754), .b(n1750), .O(n1755));
  orx  g1715(.a(n1755), .b(n244), .O(n1756));
  andx g1716(.a(n1454), .b(n120), .O(n1757));
  andx g1717(.a(n1687), .b(n63), .O(n1758));
  andx g1718(.a(n1695), .b(n67), .O(n1759));
  andx g1719(.a(n1759), .b(n1758), .O(n1760));
  andx g1720(.a(n1760), .b(n1757), .O(n1761));
  andx g1721(.a(n278), .b(n44), .O(n1762));
  andx g1722(.a(n1694), .b(n119), .O(n1763));
  andx g1723(.a(n1763), .b(n1762), .O(n1764));
  andx g1724(.a(n1764), .b(n1761), .O(n1765));
  andx g1725(.a(pi37), .b(n303), .O(n1766));
  andx g1726(.a(n1766), .b(n139), .O(n1767));
  andx g1727(.a(n93), .b(n91), .O(n1768));
  andx g1728(.a(n1768), .b(n278), .O(n1769));
  andx g1729(.a(n1769), .b(n1767), .O(n1770));
  andx g1730(.a(n1695), .b(n66), .O(n1771));
  andx g1731(.a(n1771), .b(n59), .O(n1772));
  andx g1732(.a(n88), .b(n1687), .O(n1773));
  andx g1733(.a(n1773), .b(n229), .O(n1774));
  andx g1734(.a(n1774), .b(n1772), .O(n1775));
  andx g1735(.a(n1775), .b(n1770), .O(n1776));
  orx  g1736(.a(n1776), .b(n1765), .O(n1777));
  andx g1737(.a(n313), .b(n307), .O(n1778));
  andx g1738(.a(n1778), .b(n254), .O(n1779));
  andx g1739(.a(pi37), .b(n63), .O(n1780));
  andx g1740(.a(n1780), .b(n66), .O(n1781));
  andx g1741(.a(n345), .b(n328), .O(n1782));
  andx g1742(.a(n1782), .b(n1781), .O(n1783));
  andx g1743(.a(n1783), .b(n1779), .O(n1784));
  andx g1744(.a(n1544), .b(n72), .O(n1785));
  andx g1745(.a(pi37), .b(n67), .O(n1786));
  andx g1746(.a(n80), .b(n64), .O(n1787));
  andx g1747(.a(n1787), .b(n1786), .O(n1788));
  andx g1748(.a(n351), .b(n147), .O(n1789));
  andx g1749(.a(n1789), .b(n1788), .O(n1790));
  andx g1750(.a(n1790), .b(n1785), .O(n1791));
  orx  g1751(.a(n1791), .b(n1784), .O(n1792));
  orx  g1752(.a(n1792), .b(n1777), .O(n1793));
  orx  g1753(.a(n1793), .b(n1756), .O(n1794));
  andx g1754(.a(n1344), .b(n117), .O(n1795));
  andx g1755(.a(pi10), .b(n63), .O(n1796));
  andx g1756(.a(n1796), .b(n1753), .O(n1797));
  andx g1757(.a(n1797), .b(n130), .O(n1798));
  andx g1758(.a(n1798), .b(n1795), .O(n1799));
  orx  g1759(.a(n1799), .b(n354), .O(n1800));
  andx g1760(.a(pi27), .b(n57), .O(n1801));
  andx g1761(.a(n80), .b(n56), .O(n1802));
  andx g1762(.a(n1802), .b(n1801), .O(n1803));
  andx g1763(.a(n248), .b(n90), .O(n1804));
  andx g1764(.a(n1804), .b(n1803), .O(n1805));
  andx g1765(.a(n1805), .b(n200), .O(n1806));
  orx  g1766(.a(n1806), .b(n1283), .O(n1807));
  orx  g1767(.a(n1807), .b(n1800), .O(n1808));
  andx g1768(.a(n1751), .b(n1039), .O(n1809));
  andx g1769(.a(n65), .b(n87), .O(n1810));
  andx g1770(.a(pi37), .b(n1687), .O(n1811));
  andx g1771(.a(n1811), .b(n1610), .O(n1812));
  andx g1772(.a(n1812), .b(n1810), .O(n1813));
  andx g1773(.a(n1813), .b(n1809), .O(n1814));
  andx g1774(.a(pi09), .b(pi11), .O(n1815));
  andx g1775(.a(n1815), .b(n207), .O(n1816));
  andx g1776(.a(n1816), .b(n1198), .O(n1817));
  andx g1777(.a(n1786), .b(n238), .O(n1818));
  andx g1778(.a(n1818), .b(n712), .O(n1819));
  andx g1779(.a(n1819), .b(n1817), .O(n1820));
  orx  g1780(.a(n1820), .b(n1814), .O(n1821));
  orx  g1781(.a(n1821), .b(n1313), .O(n1822));
  orx  g1782(.a(n1822), .b(n1808), .O(n1823));
  orx  g1783(.a(n1823), .b(n1794), .O(n1824));
  orx  g1784(.a(n1824), .b(n1747), .O(n1825));
  andx g1785(.a(n943), .b(n42), .O(n1826));
  andx g1786(.a(n1826), .b(n52), .O(n1827));
  andx g1787(.a(pi09), .b(n57), .O(n1828));
  andx g1788(.a(n1828), .b(n127), .O(n1829));
  andx g1789(.a(n1758), .b(n61), .O(n1830));
  andx g1790(.a(n533), .b(n64), .O(n1831));
  andx g1791(.a(pi37), .b(n66), .O(n1832));
  andx g1792(.a(n1832), .b(n1831), .O(n1833));
  andx g1793(.a(n1833), .b(n1830), .O(n1834));
  andx g1794(.a(n1834), .b(n1829), .O(n1835));
  andx g1795(.a(n1835), .b(n1827), .O(n1836));
  andx g1796(.a(n1826), .b(pi07), .O(n1837));
  andx g1797(.a(pi37), .b(n64), .O(n1838));
  andx g1798(.a(n1838), .b(n749), .O(n1839));
  andx g1799(.a(n1839), .b(n292), .O(n1840));
  andx g1800(.a(n1840), .b(n108), .O(n1841));
  andx g1801(.a(n1841), .b(n1837), .O(n1842));
  orx  g1802(.a(n1842), .b(n1836), .O(n1843));
  andx g1803(.a(n49), .b(n1695), .O(n1844));
  andx g1804(.a(n1844), .b(pi29), .O(n1845));
  andx g1805(.a(n1845), .b(pi37), .O(n1846));
  andx g1806(.a(n935), .b(n107), .O(n1847));
  andx g1807(.a(n214), .b(n277), .O(n1848));
  andx g1808(.a(n1848), .b(n117), .O(n1849));
  andx g1809(.a(n1849), .b(n1847), .O(n1850));
  andx g1810(.a(n450), .b(n264), .O(n1851));
  andx g1811(.a(n1851), .b(n1850), .O(n1852));
  andx g1812(.a(n1852), .b(n1846), .O(n1853));
  andx g1813(.a(n1811), .b(n119), .O(n1854));
  andx g1814(.a(n1831), .b(n229), .O(n1855));
  andx g1815(.a(n1855), .b(n1854), .O(n1856));
  andx g1816(.a(n1856), .b(n807), .O(n1857));
  andx g1817(.a(n1857), .b(n1837), .O(n1858));
  orx  g1818(.a(n1858), .b(n1853), .O(n1859));
  orx  g1819(.a(n1859), .b(n1843), .O(n1860));
  andx g1820(.a(n229), .b(n207), .O(n1861));
  andx g1821(.a(n1710), .b(n369), .O(n1862));
  andx g1822(.a(n1862), .b(n1861), .O(n1863));
  andx g1823(.a(n1863), .b(n1712), .O(n1864));
  andx g1824(.a(n240), .b(n182), .O(n1865));
  andx g1825(.a(n1865), .b(n1732), .O(n1866));
  andx g1826(.a(n1866), .b(n1731), .O(n1867));
  orx  g1827(.a(n1867), .b(n1864), .O(n1868));
  andx g1828(.a(n895), .b(n144), .O(n1869));
  andx g1829(.a(n277), .b(n57), .O(n1870));
  andx g1830(.a(n1870), .b(n1454), .O(n1871));
  andx g1831(.a(n1871), .b(n1869), .O(n1872));
  andx g1832(.a(n1305), .b(n1697), .O(n1873));
  andx g1833(.a(n1873), .b(n1872), .O(n1874));
  orx  g1834(.a(n1874), .b(n1402), .O(n1875));
  orx  g1835(.a(n1875), .b(n1868), .O(n1876));
  andx g1836(.a(n89), .b(n52), .O(n1877));
  andx g1837(.a(n1877), .b(n584), .O(n1878));
  andx g1838(.a(n1878), .b(n994), .O(n1879));
  orx  g1839(.a(n1879), .b(n1522), .O(n1880));
  andx g1840(.a(n1344), .b(n220), .O(n1881));
  andx g1841(.a(n1881), .b(n1720), .O(n1882));
  andx g1842(.a(n1882), .b(n1389), .O(n1883));
  andx g1843(.a(n59), .b(pi27), .O(n1884));
  andx g1844(.a(n1884), .b(n58), .O(n1885));
  andx g1845(.a(n1885), .b(n1725), .O(n1886));
  andx g1846(.a(n200), .b(n204), .O(n1887));
  andx g1847(.a(n1887), .b(n1886), .O(n1888));
  orx  g1848(.a(n1888), .b(n1883), .O(n1889));
  orx  g1849(.a(n1889), .b(n1880), .O(n1890));
  orx  g1850(.a(n1890), .b(n1876), .O(n1891));
  andx g1851(.a(n1795), .b(n60), .O(n1892));
  andx g1852(.a(n1753), .b(n63), .O(n1893));
  andx g1853(.a(n1893), .b(n248), .O(n1894));
  andx g1854(.a(n1894), .b(n1892), .O(n1895));
  andx g1855(.a(n653), .b(n345), .O(n1896));
  andx g1856(.a(n1896), .b(n1752), .O(n1897));
  andx g1857(.a(n1838), .b(n76), .O(n1898));
  andx g1858(.a(n1898), .b(n1344), .O(n1899));
  andx g1859(.a(n1802), .b(n63), .O(n1900));
  andx g1860(.a(n67), .b(n91), .O(n1901));
  andx g1861(.a(n1901), .b(n694), .O(n1902));
  andx g1862(.a(n1902), .b(n1900), .O(n1903));
  andx g1863(.a(n1903), .b(n1899), .O(n1904));
  orx  g1864(.a(n1904), .b(n1897), .O(n1905));
  orx  g1865(.a(n1905), .b(n1895), .O(n1906));
  andx g1866(.a(n163), .b(pi27), .O(n1907));
  andx g1867(.a(n238), .b(n63), .O(n1908));
  andx g1868(.a(pi10), .b(pi09), .O(n1909));
  andx g1869(.a(n1909), .b(n147), .O(n1910));
  andx g1870(.a(n1910), .b(n1908), .O(n1911));
  andx g1871(.a(n1911), .b(n1907), .O(n1912));
  andx g1872(.a(n238), .b(n64), .O(n1913));
  andx g1873(.a(n1913), .b(n1910), .O(n1914));
  andx g1874(.a(n1914), .b(n189), .O(n1915));
  orx  g1875(.a(n1915), .b(n1912), .O(n1916));
  andx g1876(.a(n60), .b(n88), .O(n1917));
  andx g1877(.a(n1917), .b(n248), .O(n1918));
  andx g1878(.a(n1918), .b(n200), .O(n1919));
  andx g1879(.a(n1919), .b(n1907), .O(n1920));
  andx g1880(.a(pi37), .b(n56), .O(n1921));
  andx g1881(.a(n1921), .b(n92), .O(n1922));
  andx g1882(.a(n1922), .b(n1870), .O(n1923));
  andx g1883(.a(n1759), .b(n432), .O(n1924));
  andx g1884(.a(n1924), .b(n1191), .O(n1925));
  andx g1885(.a(n1925), .b(n1923), .O(n1926));
  orx  g1886(.a(n1926), .b(n1920), .O(n1927));
  orx  g1887(.a(n1927), .b(n1916), .O(n1928));
  orx  g1888(.a(n1928), .b(n1906), .O(n1929));
  orx  g1889(.a(n1929), .b(n1891), .O(n1930));
  orx  g1890(.a(n1930), .b(n1860), .O(n1931));
  orx  g1891(.a(n1931), .b(n1825), .O(n1932));
  andx g1892(.a(n995), .b(n257), .O(n1933));
  andx g1893(.a(n240), .b(n171), .O(n1934));
  andx g1894(.a(n1934), .b(n1933), .O(n1935));
  andx g1895(.a(n1935), .b(n1900), .O(n1936));
  orx  g1896(.a(n1936), .b(n261), .O(n1937));
  andx g1897(.a(n1884), .b(n1725), .O(n1938));
  andx g1898(.a(n1938), .b(n375), .O(n1939));
  andx g1899(.a(n1706), .b(n171), .O(n1940));
  andx g1900(.a(n1940), .b(n1939), .O(n1941));
  andx g1901(.a(n67), .b(n63), .O(n1942));
  andx g1902(.a(n1942), .b(n1838), .O(n1943));
  andx g1903(.a(n351), .b(n130), .O(n1944));
  andx g1904(.a(n1944), .b(n1943), .O(n1945));
  andx g1905(.a(n1945), .b(n1705), .O(n1946));
  orx  g1906(.a(n1946), .b(n1941), .O(n1947));
  orx  g1907(.a(n1947), .b(n1937), .O(n1948));
  andx g1908(.a(n430), .b(n351), .O(n1949));
  andx g1909(.a(n1949), .b(n484), .O(n1950));
  andx g1910(.a(n171), .b(n117), .O(n1951));
  andx g1911(.a(n1780), .b(n80), .O(n1952));
  andx g1912(.a(n1952), .b(n1951), .O(n1953));
  andx g1913(.a(n1953), .b(n1950), .O(n1954));
  andx g1914(.a(n269), .b(pi37), .O(n1955));
  andx g1915(.a(n895), .b(n229), .O(n1956));
  andx g1916(.a(n1688), .b(n557), .O(n1957));
  andx g1917(.a(n1957), .b(n1956), .O(n1958));
  andx g1918(.a(n1958), .b(n1955), .O(n1959));
  orx  g1919(.a(n1959), .b(n1954), .O(n1960));
  orx  g1920(.a(n1960), .b(n372), .O(n1961));
  orx  g1921(.a(n1961), .b(n1948), .O(n1962));
  andx g1922(.a(n1780), .b(n345), .O(n1963));
  andx g1923(.a(n1963), .b(n392), .O(n1964));
  andx g1924(.a(n1964), .b(n96), .O(n1965));
  andx g1925(.a(n381), .b(n63), .O(n1966));
  andx g1926(.a(n1733), .b(n1730), .O(n1967));
  andx g1927(.a(n1967), .b(n1442), .O(n1968));
  andx g1928(.a(n1968), .b(n1966), .O(n1969));
  orx  g1929(.a(n1969), .b(n1965), .O(n1970));
  andx g1930(.a(n1786), .b(n902), .O(n1971));
  andx g1931(.a(n269), .b(n130), .O(n1972));
  andx g1932(.a(n1972), .b(n1971), .O(n1973));
  andx g1933(.a(n1973), .b(n700), .O(n1974));
  andx g1934(.a(n328), .b(n120), .O(n1975));
  andx g1935(.a(n303), .b(n277), .O(n1976));
  andx g1936(.a(n1976), .b(n1771), .O(n1977));
  andx g1937(.a(n1977), .b(n1975), .O(n1978));
  andx g1938(.a(n1780), .b(n67), .O(n1979));
  andx g1939(.a(n1979), .b(n1544), .O(n1980));
  andx g1940(.a(n1980), .b(n1978), .O(n1981));
  orx  g1941(.a(n1981), .b(n1974), .O(n1982));
  orx  g1942(.a(n1982), .b(n1970), .O(n1983));
  andx g1943(.a(n1802), .b(n995), .O(n1984));
  andx g1944(.a(n240), .b(n72), .O(n1985));
  andx g1945(.a(n1985), .b(n1984), .O(n1986));
  andx g1946(.a(n1986), .b(n1514), .O(n1987));
  andx g1947(.a(n238), .b(n91), .O(n1988));
  andx g1948(.a(n1838), .b(n895), .O(n1989));
  andx g1949(.a(n557), .b(n229), .O(n1990));
  andx g1950(.a(n1990), .b(n1989), .O(n1991));
  andx g1951(.a(n1991), .b(n1988), .O(n1992));
  orx  g1952(.a(n1992), .b(n1987), .O(n1993));
  andx g1953(.a(n345), .b(n248), .O(n1994));
  andx g1954(.a(n1994), .b(n53), .O(n1995));
  andx g1955(.a(n1995), .b(n190), .O(n1996));
  andx g1956(.a(n254), .b(n57), .O(n1997));
  andx g1957(.a(n274), .b(n228), .O(n1998));
  andx g1958(.a(n277), .b(n63), .O(n1999));
  andx g1959(.a(n1999), .b(n1802), .O(n2000));
  andx g1960(.a(n2000), .b(n1998), .O(n2001));
  andx g1961(.a(n2001), .b(n1997), .O(n2002));
  orx  g1962(.a(n2002), .b(n1996), .O(n2003));
  orx  g1963(.a(n2003), .b(n1993), .O(n2004));
  orx  g1964(.a(n2004), .b(n1983), .O(n2005));
  orx  g1965(.a(n2005), .b(n1962), .O(n2006));
  andx g1966(.a(n449), .b(n351), .O(n2007));
  andx g1967(.a(n2007), .b(n1811), .O(n2008));
  andx g1968(.a(n2008), .b(n105), .O(n2009));
  andx g1969(.a(n2009), .b(n1362), .O(n2010));
  andx g1970(.a(n1844), .b(n67), .O(n2011));
  andx g1971(.a(n533), .b(n59), .O(n2012));
  andx g1972(.a(n2012), .b(n268), .O(n2013));
  andx g1973(.a(n2013), .b(n1832), .O(n2014));
  andx g1974(.a(n1870), .b(n107), .O(n2015));
  andx g1975(.a(n75), .b(n56), .O(n2016));
  andx g1976(.a(n2016), .b(n491), .O(n2017));
  andx g1977(.a(n2017), .b(n2015), .O(n2018));
  andx g1978(.a(n2018), .b(n2014), .O(n2019));
  andx g1979(.a(n2019), .b(n2011), .O(n2020));
  orx  g1980(.a(n2020), .b(n2010), .O(n2021));
  andx g1981(.a(n88), .b(n91), .O(n2022));
  andx g1982(.a(n2022), .b(n315), .O(n2023));
  andx g1983(.a(n171), .b(n64), .O(n2024));
  andx g1984(.a(n1811), .b(n1706), .O(n2025));
  andx g1985(.a(n2025), .b(n2024), .O(n2026));
  andx g1986(.a(n2026), .b(n2023), .O(n2027));
  andx g1987(.a(n1844), .b(pi37), .O(n2028));
  andx g1988(.a(n2012), .b(n1519), .O(n2029));
  andx g1989(.a(n57), .b(n87), .O(n2030));
  andx g1990(.a(n2030), .b(n93), .O(n2031));
  andx g1991(.a(n75), .b(n277), .O(n2032));
  andx g1992(.a(n2032), .b(n127), .O(n2033));
  andx g1993(.a(n2033), .b(n2031), .O(n2034));
  andx g1994(.a(n2034), .b(n2029), .O(n2035));
  andx g1995(.a(n2035), .b(n2028), .O(n2036));
  orx  g1996(.a(n2036), .b(n2027), .O(n2037));
  orx  g1997(.a(n2037), .b(n2021), .O(n2038));
  andx g1998(.a(n299), .b(n1695), .O(n2039));
  andx g1999(.a(n2039), .b(n303), .O(n2040));
  andx g2000(.a(n2040), .b(n2019), .O(n2041));
  andx g2001(.a(n250), .b(n245), .O(n2042));
  andx g2002(.a(n268), .b(n53), .O(n2043));
  andx g2003(.a(n2043), .b(n2042), .O(n2044));
  andx g2004(.a(n59), .b(n277), .O(n2045));
  andx g2005(.a(n2045), .b(n58), .O(n2046));
  andx g2006(.a(n369), .b(n274), .O(n2047));
  andx g2007(.a(n2047), .b(n286), .O(n2048));
  andx g2008(.a(n2048), .b(n2046), .O(n2049));
  orx  g2009(.a(n2049), .b(n2044), .O(n2050));
  orx  g2010(.a(n2050), .b(n2041), .O(n2051));
  andx g2011(.a(n1688), .b(n53), .O(n2052));
  andx g2012(.a(n2052), .b(n1781), .O(n2053));
  andx g2013(.a(n2053), .b(n2023), .O(n2054));
  andx g2014(.a(n1811), .b(n1198), .O(n2055));
  andx g2015(.a(n2055), .b(n53), .O(n2056));
  andx g2016(.a(n2056), .b(n712), .O(n2057));
  andx g2017(.a(n2057), .b(n1362), .O(n2058));
  orx  g2018(.a(n2058), .b(n2054), .O(n2059));
  orx  g2019(.a(n2059), .b(n2051), .O(n2060));
  orx  g2020(.a(n2060), .b(n2038), .O(n2061));
  orx  g2021(.a(n2061), .b(n2006), .O(n2062));
  andx g2022(.a(n60), .b(pi23), .O(n2063));
  andx g2023(.a(n2063), .b(n1885), .O(n2064));
  andx g2024(.a(n286), .b(n257), .O(n2065));
  andx g2025(.a(n2065), .b(n2064), .O(n2066));
  andx g2026(.a(n1832), .b(n1759), .O(n2067));
  andx g2027(.a(n2067), .b(n2045), .O(n2068));
  andx g2028(.a(n491), .b(n92), .O(n2069));
  andx g2029(.a(n2069), .b(n1861), .O(n2070));
  andx g2030(.a(n2070), .b(n2068), .O(n2071));
  orx  g2031(.a(n2071), .b(n2066), .O(n2072));
  andx g2032(.a(n1766), .b(n207), .O(n2073));
  andx g2033(.a(n2045), .b(n1503), .O(n2074));
  andx g2034(.a(n2074), .b(n2073), .O(n2075));
  andx g2035(.a(n1758), .b(n75), .O(n2076));
  andx g2036(.a(n1759), .b(n119), .O(n2077));
  andx g2037(.a(n2077), .b(n2076), .O(n2078));
  andx g2038(.a(n2078), .b(n2075), .O(n2079));
  andx g2039(.a(n1951), .b(n60), .O(n2080));
  andx g2040(.a(n1740), .b(n63), .O(n2081));
  andx g2041(.a(n2081), .b(n125), .O(n2082));
  andx g2042(.a(n2082), .b(n2080), .O(n2083));
  orx  g2043(.a(n2083), .b(n2079), .O(n2084));
  orx  g2044(.a(n2084), .b(n2072), .O(n2085));
  andx g2045(.a(n1710), .b(n273), .O(n2086));
  andx g2046(.a(n2086), .b(n1861), .O(n2087));
  andx g2047(.a(n2087), .b(n1712), .O(n2088));
  andx g2048(.a(n1544), .b(pi27), .O(n2089));
  andx g2049(.a(n204), .b(pi07), .O(n2090));
  andx g2050(.a(n1796), .b(n147), .O(n2091));
  andx g2051(.a(n2091), .b(n2090), .O(n2092));
  andx g2052(.a(n2092), .b(n2089), .O(n2093));
  orx  g2053(.a(n2093), .b(n2088), .O(n2094));
  andx g2054(.a(n171), .b(n59), .O(n2095));
  andx g2055(.a(n268), .b(n139), .O(n2096));
  andx g2056(.a(n2096), .b(n2095), .O(n2097));
  andx g2057(.a(n2097), .b(n1711), .O(n2098));
  orx  g2058(.a(n2098), .b(n1373), .O(n2099));
  orx  g2059(.a(n2099), .b(n2094), .O(n2100));
  orx  g2060(.a(n2100), .b(n2085), .O(n2101));
  andx g2061(.a(n397), .b(n66), .O(n2102));
  andx g2062(.a(n2102), .b(n182), .O(n2103));
  andx g2063(.a(n2103), .b(n1886), .O(n2104));
  orx  g2064(.a(n2104), .b(n1391), .O(n2105));
  andx g2065(.a(n1454), .b(n491), .O(n2106));
  andx g2066(.a(n1780), .b(n484), .O(n2107));
  andx g2067(.a(n2107), .b(n2106), .O(n2108));
  andx g2068(.a(n1772), .b(n1762), .O(n2109));
  andx g2069(.a(n2109), .b(n2108), .O(n2110));
  orx  g2070(.a(n2110), .b(n288), .O(n2111));
  orx  g2071(.a(n2111), .b(n2105), .O(n2112));
  andx g2072(.a(n855), .b(n328), .O(n2113));
  andx g2073(.a(n2113), .b(n484), .O(n2114));
  andx g2074(.a(n1838), .b(n66), .O(n2115));
  andx g2075(.a(n2115), .b(n1795), .O(n2116));
  andx g2076(.a(n2116), .b(n2114), .O(n2117));
  andx g2077(.a(n1766), .b(n1688), .O(n2118));
  andx g2078(.a(n2118), .b(n653), .O(n2119));
  andx g2079(.a(n2119), .b(n1809), .O(n2120));
  orx  g2080(.a(n2120), .b(n2117), .O(n2121));
  andx g2081(.a(n248), .b(n204), .O(n2122));
  andx g2082(.a(n1392), .b(n323), .O(n2123));
  andx g2083(.a(n2123), .b(n2122), .O(n2124));
  andx g2084(.a(n2124), .b(n1997), .O(n2125));
  andx g2085(.a(pi37), .b(n249), .O(n2126));
  andx g2086(.a(n2126), .b(n53), .O(n2127));
  andx g2087(.a(n164), .b(n92), .O(n2128));
  andx g2088(.a(n2128), .b(n397), .O(n2129));
  andx g2089(.a(n2129), .b(n2127), .O(n2130));
  orx  g2090(.a(n2130), .b(n2125), .O(n2131));
  orx  g2091(.a(n2131), .b(n2121), .O(n2132));
  orx  g2092(.a(n2132), .b(n2112), .O(n2133));
  orx  g2093(.a(n2133), .b(n2101), .O(n2134));
  andx g2094(.a(n80), .b(pi07), .O(n2135));
  andx g2095(.a(n2135), .b(n64), .O(n2136));
  andx g2096(.a(n2136), .b(n2091), .O(n2137));
  andx g2097(.a(n2137), .b(n1951), .O(n2138));
  orx  g2098(.a(n2138), .b(n1516), .O(n2139));
  andx g2099(.a(n1921), .b(n1768), .O(n2140));
  andx g2100(.a(n2140), .b(n1870), .O(n2141));
  andx g2101(.a(n1204), .b(n431), .O(n2142));
  andx g2102(.a(n1771), .b(n432), .O(n2143));
  andx g2103(.a(n2143), .b(n2142), .O(n2144));
  andx g2104(.a(n2144), .b(n2141), .O(n2145));
  orx  g2105(.a(n2145), .b(n1531), .O(n2146));
  orx  g2106(.a(n2146), .b(n2139), .O(n2147));
  andx g2107(.a(n1725), .b(n144), .O(n2148));
  andx g2108(.a(n2148), .b(n1801), .O(n2149));
  andx g2109(.a(pi09), .b(n59), .O(n2150));
  andx g2110(.a(n2150), .b(n690), .O(n2151));
  andx g2111(.a(n2151), .b(n2149), .O(n2152));
  andx g2112(.a(n1280), .b(n200), .O(n2153));
  andx g2113(.a(n2153), .b(n2064), .O(n2154));
  orx  g2114(.a(n2154), .b(n2152), .O(n2155));
  andx g2115(.a(n286), .b(n206), .O(n2156));
  andx g2116(.a(n2156), .b(n2149), .O(n2157));
  andx g2117(.a(n1706), .b(n345), .O(n2158));
  andx g2118(.a(n2158), .b(n248), .O(n2159));
  andx g2119(.a(n2159), .b(n2080), .O(n2160));
  orx  g2120(.a(n2160), .b(n2157), .O(n2161));
  orx  g2121(.a(n2161), .b(n2155), .O(n2162));
  orx  g2122(.a(n2162), .b(n2147), .O(n2163));
  andx g2123(.a(n72), .b(n53), .O(n2164));
  andx g2124(.a(n2164), .b(n1939), .O(n2165));
  andx g2125(.a(n432), .b(n67), .O(n2166));
  andx g2126(.a(n545), .b(n104), .O(n2167));
  andx g2127(.a(n1838), .b(n250), .O(n2168));
  andx g2128(.a(n2168), .b(n2167), .O(n2169));
  andx g2129(.a(n2169), .b(n2166), .O(n2170));
  orx  g2130(.a(n2170), .b(n2165), .O(n2171));
  andx g2131(.a(n1918), .b(n653), .O(n2172));
  andx g2132(.a(n2172), .b(n2089), .O(n2173));
  andx g2133(.a(n1740), .b(n80), .O(n2174));
  andx g2134(.a(n2174), .b(n125), .O(n2175));
  andx g2135(.a(n2175), .b(n1785), .O(n2176));
  orx  g2136(.a(n2176), .b(n2173), .O(n2177));
  orx  g2137(.a(n2177), .b(n2171), .O(n2178));
  andx g2138(.a(n1768), .b(n1766), .O(n2179));
  andx g2139(.a(n2179), .b(n2045), .O(n2180));
  andx g2140(.a(n1771), .b(n491), .O(n2181));
  andx g2141(.a(n2181), .b(n1861), .O(n2182));
  andx g2142(.a(n2182), .b(n2180), .O(n2183));
  andx g2143(.a(n1771), .b(n328), .O(n2184));
  andx g2144(.a(n2184), .b(n895), .O(n2185));
  andx g2145(.a(n1780), .b(n1344), .O(n2186));
  andx g2146(.a(n2186), .b(n2046), .O(n2187));
  andx g2147(.a(n2187), .b(n2185), .O(n2188));
  orx  g2148(.a(n2188), .b(n2183), .O(n2189));
  andx g2149(.a(n1344), .b(n207), .O(n2190));
  andx g2150(.a(n2190), .b(n589), .O(n2191));
  andx g2151(.a(n1198), .b(n130), .O(n2192));
  andx g2152(.a(n2192), .b(n1979), .O(n2193));
  andx g2153(.a(n2193), .b(n2191), .O(n2194));
  andx g2154(.a(n1786), .b(n199), .O(n2195));
  andx g2155(.a(n52), .b(n249), .O(n2196));
  andx g2156(.a(n1688), .b(n92), .O(n2197));
  andx g2157(.a(n2197), .b(n2196), .O(n2198));
  andx g2158(.a(n2198), .b(n2195), .O(n2199));
  orx  g2159(.a(n2199), .b(n2194), .O(n2200));
  orx  g2160(.a(n2200), .b(n2189), .O(n2201));
  orx  g2161(.a(n2201), .b(n2178), .O(n2202));
  orx  g2162(.a(n2202), .b(n2163), .O(n2203));
  orx  g2163(.a(n2203), .b(n2134), .O(n2204));
  orx  g2164(.a(n2204), .b(n2062), .O(n2205));
  orx  g2165(.a(n2205), .b(n1932), .O(n2206));
  andx g2166(.a(n677), .b(n42), .O(n2207));
  andx g2167(.a(n2207), .b(pi07), .O(n2208));
  andx g2168(.a(n1687), .b(n57), .O(n2209));
  andx g2169(.a(n2209), .b(n254), .O(n2210));
  andx g2170(.a(n1921), .b(n647), .O(n2211));
  andx g2171(.a(n2211), .b(n69), .O(n2212));
  andx g2172(.a(n2212), .b(n2210), .O(n2213));
  andx g2173(.a(n2213), .b(n2208), .O(n2214));
  andx g2174(.a(n813), .b(n1695), .O(n2215));
  andx g2175(.a(n2215), .b(pi37), .O(n2216));
  andx g2176(.a(n2216), .b(n895), .O(n2217));
  andx g2177(.a(n1999), .b(n76), .O(n2218));
  andx g2178(.a(n1687), .b(n56), .O(n2219));
  andx g2179(.a(n2219), .b(n1080), .O(n2220));
  andx g2180(.a(n647), .b(n171), .O(n2221));
  andx g2181(.a(n2221), .b(n2220), .O(n2222));
  andx g2182(.a(n2222), .b(n2218), .O(n2223));
  andx g2183(.a(n2223), .b(n2217), .O(n2224));
  orx  g2184(.a(n2224), .b(n2214), .O(n2225));
  andx g2185(.a(n1828), .b(n107), .O(n2226));
  andx g2186(.a(n1921), .b(n65), .O(n2227));
  andx g2187(.a(n2227), .b(n984), .O(n2228));
  andx g2188(.a(n2228), .b(n2226), .O(n2229));
  andx g2189(.a(n2229), .b(n1827), .O(n2230));
  andx g2190(.a(n80), .b(n42), .O(n2231));
  andx g2191(.a(n730), .b(n303), .O(n2232));
  andx g2192(.a(n2232), .b(n2231), .O(n2233));
  andx g2193(.a(n733), .b(n87), .O(n2234));
  andx g2194(.a(n735), .b(n449), .O(n2235));
  andx g2195(.a(n1694), .b(n494), .O(n2236));
  andx g2196(.a(n2236), .b(n2235), .O(n2237));
  andx g2197(.a(n2237), .b(n2234), .O(n2238));
  andx g2198(.a(n2238), .b(n2233), .O(n2239));
  orx  g2199(.a(n2239), .b(n2230), .O(n2240));
  orx  g2200(.a(n2240), .b(n2225), .O(n2241));
  andx g2201(.a(n2207), .b(n52), .O(n2242));
  andx g2202(.a(n1921), .b(n1758), .O(n2243));
  andx g2203(.a(n1831), .b(n381), .O(n2244));
  andx g2204(.a(n2244), .b(n2243), .O(n2245));
  andx g2205(.a(n2245), .b(n624), .O(n2246));
  andx g2206(.a(n2246), .b(n2242), .O(n2247));
  andx g2207(.a(n2231), .b(n677), .O(n2248));
  andx g2208(.a(n2248), .b(pi07), .O(n2249));
  andx g2209(.a(n117), .b(n68), .O(n2250));
  andx g2210(.a(n1838), .b(n229), .O(n2251));
  andx g2211(.a(n2251), .b(n2250), .O(n2252));
  andx g2212(.a(n2252), .b(n1211), .O(n2253));
  andx g2213(.a(n2253), .b(n2249), .O(n2254));
  orx  g2214(.a(n2254), .b(n2247), .O(n2255));
  andx g2215(.a(n214), .b(n212), .O(n2256));
  andx g2216(.a(n2256), .b(n1870), .O(n2257));
  andx g2217(.a(n59), .b(n87), .O(n2258));
  andx g2218(.a(n2258), .b(n204), .O(n2259));
  andx g2219(.a(n2016), .b(n268), .O(n2260));
  andx g2220(.a(n2260), .b(n2259), .O(n2261));
  andx g2221(.a(n2261), .b(n2257), .O(n2262));
  andx g2222(.a(n2262), .b(n2217), .O(n2263));
  andx g2223(.a(n2665), .b(n60), .O(n2264));
  andx g2224(.a(pi11), .b(n91), .O(n2265));
  andx g2225(.a(n2265), .b(n2264), .O(n2266));
  andx g2226(.a(n1786), .b(n1688), .O(n2267));
  andx g2227(.a(n2267), .b(n653), .O(n2268));
  andx g2228(.a(n2268), .b(n2266), .O(n2269));
  orx  g2229(.a(n2269), .b(n2263), .O(n2270));
  orx  g2230(.a(n2270), .b(n2255), .O(n2271));
  orx  g2231(.a(n2271), .b(n2241), .O(n2272));
  andx g2232(.a(n2231), .b(n943), .O(n2273));
  andx g2233(.a(n2273), .b(n52), .O(n2274));
  andx g2234(.a(n199), .b(n90), .O(n2275));
  andx g2235(.a(n1921), .b(n345), .O(n2276));
  andx g2236(.a(n2276), .b(n2275), .O(n2277));
  andx g2237(.a(n2277), .b(n2274), .O(n2278));
  andx g2238(.a(n730), .b(n42), .O(n2279));
  andx g2239(.a(n2279), .b(pi07), .O(n2280));
  andx g2240(.a(n76), .b(pi26), .O(n2281));
  andx g2241(.a(n449), .b(n397), .O(n2282));
  andx g2242(.a(n1921), .b(n1610), .O(n2283));
  andx g2243(.a(n2283), .b(n2282), .O(n2284));
  andx g2244(.a(n2284), .b(n2281), .O(n2285));
  andx g2245(.a(n2285), .b(n2280), .O(n2286));
  orx  g2246(.a(n2286), .b(n2278), .O(n2287));
  andx g2247(.a(n494), .b(n107), .O(n2288));
  andx g2248(.a(n1921), .b(n589), .O(n2289));
  andx g2249(.a(n2289), .b(n1124), .O(n2290));
  andx g2250(.a(n2290), .b(n2288), .O(n2291));
  andx g2251(.a(n2291), .b(n2274), .O(n2292));
  andx g2252(.a(n1802), .b(n229), .O(n2293));
  andx g2253(.a(n1832), .b(n164), .O(n2294));
  andx g2254(.a(n2294), .b(n2293), .O(n2295));
  andx g2255(.a(n2295), .b(n2281), .O(n2296));
  andx g2256(.a(n2296), .b(n2208), .O(n2297));
  orx  g2257(.a(n2297), .b(n2292), .O(n2298));
  orx  g2258(.a(n2298), .b(n2287), .O(n2299));
  andx g2259(.a(n60), .b(n277), .O(n2300));
  andx g2260(.a(n2300), .b(n2030), .O(n2301));
  andx g2261(.a(n1758), .b(n117), .O(n2302));
  andx g2262(.a(n41), .b(pi29), .O(n2303));
  andx g2263(.a(n2303), .b(n171), .O(n2304));
  andx g2264(.a(n2304), .b(n2302), .O(n2305));
  andx g2265(.a(n2305), .b(n2301), .O(n2306));
  andx g2266(.a(n2028), .b(n67), .O(n2307));
  andx g2267(.a(n2307), .b(n2306), .O(n2308));
  andx g2268(.a(n2231), .b(n730), .O(n2309));
  andx g2269(.a(n2309), .b(pi07), .O(n2310));
  andx g2270(.a(n171), .b(n56), .O(n2311));
  andx g2271(.a(n1780), .b(n1148), .O(n2312));
  andx g2272(.a(n2312), .b(n1667), .O(n2313));
  andx g2273(.a(n2313), .b(n2311), .O(n2314));
  andx g2274(.a(n2314), .b(n2310), .O(n2315));
  orx  g2275(.a(n2315), .b(n2308), .O(n2316));
  andx g2276(.a(n58), .b(pi26), .O(n2317));
  andx g2277(.a(n589), .b(n204), .O(n2318));
  andx g2278(.a(n2318), .b(n2195), .O(n2319));
  andx g2279(.a(n2319), .b(n2317), .O(n2320));
  andx g2280(.a(n2320), .b(n2242), .O(n2321));
  andx g2281(.a(n1205), .b(n2251), .O(n2322));
  andx g2282(.a(n2322), .b(n1211), .O(n2323));
  andx g2283(.a(n2323), .b(n2310), .O(n2324));
  orx  g2284(.a(n2324), .b(n2321), .O(n2325));
  orx  g2285(.a(n2325), .b(n2316), .O(n2326));
  orx  g2286(.a(n2326), .b(n2299), .O(n2327));
  orx  g2287(.a(n2327), .b(n2272), .O(n2328));
  andx g2288(.a(n2264), .b(pi23), .O(n2329));
  andx g2289(.a(n1280), .b(n431), .O(n2330));
  andx g2290(.a(n2330), .b(n2329), .O(n2331));
  andx g2291(.a(n421), .b(n94), .O(n2332));
  andx g2292(.a(n107), .b(n59), .O(n2333));
  andx g2293(.a(n2333), .b(n72), .O(n2334));
  andx g2294(.a(n2032), .b(n491), .O(n2335));
  andx g2295(.a(n2335), .b(n2334), .O(n2336));
  andx g2296(.a(n2336), .b(n2332), .O(n2337));
  andx g2297(.a(n2337), .b(n1846), .O(n2338));
  orx  g2298(.a(n2338), .b(n2331), .O(n2339));
  andx g2299(.a(n2016), .b(n536), .O(n2340));
  andx g2300(.a(pi26), .b(n277), .O(n2341));
  andx g2301(.a(n2341), .b(n268), .O(n2342));
  andx g2302(.a(n2342), .b(n2259), .O(n2343));
  andx g2303(.a(n2343), .b(n2340), .O(n2344));
  andx g2304(.a(n2344), .b(n2307), .O(n2345));
  andx g2305(.a(n2273), .b(pi07), .O(n2346));
  andx g2306(.a(n840), .b(n107), .O(n2347));
  andx g2307(.a(pi37), .b(n212), .O(n2348));
  andx g2308(.a(n2348), .b(n2016), .O(n2349));
  andx g2309(.a(n90), .b(n65), .O(n2350));
  andx g2310(.a(n2350), .b(n2349), .O(n2351));
  andx g2311(.a(n2351), .b(n2347), .O(n2352));
  andx g2312(.a(n2352), .b(n2346), .O(n2353));
  orx  g2313(.a(n2353), .b(n2345), .O(n2354));
  orx  g2314(.a(n2354), .b(n2339), .O(n2355));
  andx g2315(.a(n1845), .b(n1811), .O(n2356));
  andx g2316(.a(n566), .b(n72), .O(n2357));
  andx g2317(.a(n2357), .b(n2032), .O(n2358));
  andx g2318(.a(n2333), .b(n2030), .O(n2359));
  andx g2319(.a(n2359), .b(n759), .O(n2360));
  andx g2320(.a(n2360), .b(n2358), .O(n2361));
  andx g2321(.a(n2361), .b(n2356), .O(n2362));
  andx g2322(.a(n494), .b(n164), .O(n2363));
  andx g2323(.a(n1780), .b(n566), .O(n2364));
  andx g2324(.a(n2364), .b(n2363), .O(n2365));
  andx g2325(.a(n2365), .b(n1544), .O(n2366));
  andx g2326(.a(n2366), .b(n2249), .O(n2367));
  orx  g2327(.a(n2367), .b(n2362), .O(n2368));
  andx g2328(.a(n2256), .b(n428), .O(n2369));
  andx g2329(.a(n1838), .b(n104), .O(n2370));
  andx g2330(.a(n2370), .b(n2369), .O(n2371));
  andx g2331(.a(n2371), .b(n2226), .O(n2372));
  andx g2332(.a(n2372), .b(n2274), .O(n2373));
  andx g2333(.a(n1811), .b(n68), .O(n2374));
  andx g2334(.a(n2374), .b(n1810), .O(n2375));
  andx g2335(.a(n2375), .b(n2266), .O(n2376));
  orx  g2336(.a(n2376), .b(n2373), .O(n2377));
  orx  g2337(.a(n2377), .b(n2368), .O(n2378));
  orx  g2338(.a(n2378), .b(n2355), .O(n2379));
  andx g2339(.a(n2258), .b(n1921), .O(n2380));
  andx g2340(.a(n171), .b(n65), .O(n2381));
  andx g2341(.a(n2381), .b(n2380), .O(n2382));
  andx g2342(.a(n2382), .b(n1211), .O(n2383));
  andx g2343(.a(n2383), .b(n2233), .O(n2384));
  andx g2344(.a(n2248), .b(n52), .O(n2385));
  andx g2345(.a(n1828), .b(n1780), .O(n2386));
  andx g2346(.a(n566), .b(n164), .O(n2387));
  andx g2347(.a(n2387), .b(n2386), .O(n2388));
  andx g2348(.a(n2388), .b(n163), .O(n2389));
  andx g2349(.a(n2389), .b(n2385), .O(n2390));
  orx  g2350(.a(n2390), .b(n2384), .O(n2391));
  andx g2351(.a(n2030), .b(n94), .O(n2392));
  andx g2352(.a(n2032), .b(n647), .O(n2393));
  andx g2353(.a(n2393), .b(n2334), .O(n2394));
  andx g2354(.a(n2394), .b(n2392), .O(n2395));
  andx g2355(.a(n2395), .b(n2356), .O(n2396));
  andx g2356(.a(n1280), .b(n522), .O(n2397));
  andx g2357(.a(n2397), .b(n2329), .O(n2398));
  orx  g2358(.a(n2398), .b(n2396), .O(n2399));
  orx  g2359(.a(n2399), .b(n2391), .O(n2400));
  andx g2360(.a(n75), .b(n57), .O(n2401));
  andx g2361(.a(n2401), .b(n61), .O(n2402));
  andx g2362(.a(n2219), .b(n855), .O(n2403));
  andx g2363(.a(n2403), .b(n1833), .O(n2404));
  andx g2364(.a(n2404), .b(n2402), .O(n2405));
  andx g2365(.a(n2405), .b(n2280), .O(n2406));
  andx g2366(.a(n199), .b(n117), .O(n2407));
  andx g2367(.a(n2407), .b(n2294), .O(n2408));
  andx g2368(.a(n2408), .b(n1211), .O(n2409));
  andx g2369(.a(n2409), .b(n2385), .O(n2410));
  orx  g2370(.a(n2410), .b(n2406), .O(n2411));
  andx g2371(.a(n1832), .b(n254), .O(n2412));
  andx g2372(.a(n2412), .b(n208), .O(n2413));
  andx g2373(.a(n2413), .b(n2346), .O(n2414));
  andx g2374(.a(n76), .b(n107), .O(n2415));
  andx g2375(.a(n2016), .b(n566), .O(n2416));
  andx g2376(.a(n1832), .b(n65), .O(n2417));
  andx g2377(.a(n2417), .b(n2416), .O(n2418));
  andx g2378(.a(n2418), .b(n2415), .O(n2419));
  andx g2379(.a(n2419), .b(n2346), .O(n2420));
  orx  g2380(.a(n2420), .b(n2414), .O(n2421));
  orx  g2381(.a(n2421), .b(n2411), .O(n2422));
  orx  g2382(.a(n2422), .b(n2400), .O(n2423));
  orx  g2383(.a(n2423), .b(n2379), .O(n2424));
  orx  g2384(.a(n2424), .b(n2328), .O(n2425));
  orx  g2385(.a(n2425), .b(n2206), .O(n2426));
  andx g2386(.a(n891), .b(n1695), .O(n2427));
  andx g2387(.a(n277), .b(n87), .O(n2428));
  andx g2388(.a(n2428), .b(n171), .O(n2429));
  andx g2389(.a(n895), .b(n718), .O(n2430));
  andx g2390(.a(n1780), .b(n89), .O(n2431));
  andx g2391(.a(n2431), .b(n2430), .O(n2432));
  andx g2392(.a(n2432), .b(n2429), .O(n2433));
  andx g2393(.a(n2433), .b(n2427), .O(n2434));
  andx g2394(.a(n1348), .b(n41), .O(n2435));
  andx g2395(.a(n459), .b(n57), .O(n2436));
  andx g2396(.a(n2231), .b(n449), .O(n2437));
  andx g2397(.a(n1780), .b(n1204), .O(n2438));
  andx g2398(.a(n2438), .b(n2437), .O(n2439));
  andx g2399(.a(n2439), .b(n2436), .O(n2440));
  andx g2400(.a(n2440), .b(n2435), .O(n2441));
  orx  g2401(.a(n2441), .b(n2434), .O(n2442));
  andx g2402(.a(n2231), .b(n120), .O(n2443));
  andx g2403(.a(n2443), .b(n1989), .O(n2444));
  andx g2404(.a(n2444), .b(n286), .O(n2445));
  andx g2405(.a(n2445), .b(n1609), .O(n2446));
  andx g2406(.a(n1811), .b(n351), .O(n2447));
  andx g2407(.a(n2447), .b(n147), .O(n2448));
  andx g2408(.a(n2448), .b(n1343), .O(n2449));
  andx g2409(.a(n2449), .b(n2080), .O(n2450));
  orx  g2410(.a(n2450), .b(n2446), .O(n2451));
  orx  g2411(.a(n2451), .b(n2442), .O(n2452));
  andx g2412(.a(n1844), .b(n88), .O(n2453));
  andx g2413(.a(n254), .b(n87), .O(n2454));
  andx g2414(.a(n1786), .b(n228), .O(n2455));
  andx g2415(.a(n2455), .b(n2000), .O(n2456));
  andx g2416(.a(n2456), .b(n2454), .O(n2457));
  andx g2417(.a(n2457), .b(n2453), .O(n2458));
  andx g2418(.a(n943), .b(n88), .O(n2459));
  andx g2419(.a(n2219), .b(n437), .O(n2460));
  andx g2420(.a(n42), .b(pi37), .O(n2461));
  andx g2421(.a(n2461), .b(n902), .O(n2462));
  andx g2422(.a(n2462), .b(n2460), .O(n2463));
  andx g2423(.a(n2463), .b(n551), .O(n2464));
  andx g2424(.a(n2464), .b(n2459), .O(n2465));
  orx  g2425(.a(n2465), .b(n2458), .O(n2466));
  andx g2426(.a(n437), .b(n90), .O(n2467));
  andx g2427(.a(n2467), .b(n2462), .O(n2468));
  andx g2428(.a(n213), .b(n107), .O(n2469));
  andx g2429(.a(n2209), .b(n215), .O(n2470));
  andx g2430(.a(n2470), .b(n2469), .O(n2471));
  andx g2431(.a(n2471), .b(n2468), .O(n2472));
  andx g2432(.a(n2472), .b(n943), .O(n2473));
  andx g2433(.a(n1725), .b(n2665), .O(n2474));
  andx g2434(.a(n522), .b(n204), .O(n2475));
  andx g2435(.a(n2475), .b(n2474), .O(n2476));
  orx  g2436(.a(n2476), .b(n2473), .O(n2477));
  orx  g2437(.a(n2477), .b(n2466), .O(n2478));
  orx  g2438(.a(n2478), .b(n2452), .O(n2479));
  andx g2439(.a(n1666), .b(n1408), .O(n2480));
  andx g2440(.a(n1786), .b(n909), .O(n2481));
  andx g2441(.a(n2219), .b(n73), .O(n2482));
  andx g2442(.a(n2482), .b(n2481), .O(n2483));
  andx g2443(.a(n2483), .b(n2480), .O(n2484));
  andx g2444(.a(n2484), .b(n677), .O(n2485));
  andx g2445(.a(n1027), .b(n1000), .O(n2486));
  orx  g2446(.a(n2486), .b(n2485), .O(n2487));
  andx g2447(.a(n2461), .b(n2209), .O(n2488));
  andx g2448(.a(n2488), .b(n545), .O(n2489));
  andx g2449(.a(n2016), .b(n2012), .O(n2490));
  andx g2450(.a(n69), .b(n2490), .O(n2491));
  andx g2451(.a(n2491), .b(n2489), .O(n2492));
  andx g2452(.a(n2492), .b(n975), .O(n2493));
  andx g2453(.a(n2039), .b(n1811), .O(n2494));
  andx g2454(.a(n2393), .b(n108), .O(n2495));
  andx g2455(.a(n1204), .b(n72), .O(n2496));
  andx g2456(.a(n2496), .b(n1080), .O(n2497));
  andx g2457(.a(n2497), .b(n2495), .O(n2498));
  andx g2458(.a(n2498), .b(n2494), .O(n2499));
  orx  g2459(.a(n2499), .b(n2493), .O(n2500));
  orx  g2460(.a(n2500), .b(n2487), .O(n2501));
  andx g2461(.a(n1999), .b(n1766), .O(n2502));
  andx g2462(.a(n228), .b(n89), .O(n2503));
  andx g2463(.a(n2503), .b(n2502), .O(n2504));
  andx g2464(.a(n2504), .b(n1795), .O(n2505));
  andx g2465(.a(n2505), .b(n2039), .O(n2506));
  andx g2466(.a(n43), .b(n41), .O(n2507));
  andx g2467(.a(n2507), .b(n48), .O(n2508));
  andx g2468(.a(n2508), .b(n58), .O(n2509));
  andx g2469(.a(n2231), .b(n229), .O(n2510));
  andx g2470(.a(n2510), .b(n1989), .O(n2511));
  andx g2471(.a(n2511), .b(n1712), .O(n2512));
  andx g2472(.a(n2512), .b(n2509), .O(n2513));
  orx  g2473(.a(n2513), .b(n2506), .O(n2514));
  andx g2474(.a(n381), .b(n64), .O(n2515));
  andx g2475(.a(n1811), .b(n269), .O(n2516));
  andx g2476(.a(n2516), .b(n147), .O(n2517));
  andx g2477(.a(n2517), .b(n2515), .O(n2518));
  andx g2478(.a(n2518), .b(n190), .O(n2519));
  andx g2479(.a(n2231), .b(n430), .O(n2520));
  andx g2480(.a(n1780), .b(n120), .O(n2521));
  andx g2481(.a(n2521), .b(n2520), .O(n2522));
  andx g2482(.a(n2522), .b(n2095), .O(n2523));
  andx g2483(.a(n2523), .b(n1348), .O(n2524));
  orx  g2484(.a(n2524), .b(n2519), .O(n2525));
  orx  g2485(.a(n2525), .b(n2514), .O(n2526));
  orx  g2486(.a(n2526), .b(n2501), .O(n2527));
  orx  g2487(.a(n2527), .b(n2479), .O(n2528));
  andx g2488(.a(n1610), .b(n397), .O(n2529));
  andx g2489(.a(n2529), .b(n1786), .O(n2530));
  andx g2490(.a(n2341), .b(n2030), .O(n2531));
  andx g2491(.a(n404), .b(n117), .O(n2532));
  andx g2492(.a(n2532), .b(n2531), .O(n2533));
  andx g2493(.a(n2533), .b(n2530), .O(n2534));
  andx g2494(.a(n2534), .b(n2215), .O(n2535));
  andx g2495(.a(n1766), .b(n329), .O(n2536));
  andx g2496(.a(n2536), .b(n419), .O(n2537));
  andx g2497(.a(n75), .b(n212), .O(n2538));
  andx g2498(.a(n2538), .b(n2209), .O(n2539));
  andx g2499(.a(n2539), .b(n551), .O(n2540));
  andx g2500(.a(n2540), .b(n2537), .O(n2541));
  andx g2501(.a(n2541), .b(n923), .O(n2542));
  orx  g2502(.a(n2542), .b(n2535), .O(n2543));
  andx g2503(.a(n41), .b(pi07), .O(n2544));
  andx g2504(.a(n2544), .b(n2209), .O(n2545));
  andx g2505(.a(n2545), .b(n2461), .O(n2546));
  andx g2506(.a(n1213), .b(n2311), .O(n2547));
  andx g2507(.a(n2547), .b(n2546), .O(n2548));
  andx g2508(.a(n2548), .b(n1564), .O(n2549));
  andx g2509(.a(n80), .b(n41), .O(n2550));
  andx g2510(.a(n2550), .b(n1844), .O(n2551));
  andx g2511(.a(n2045), .b(n1786), .O(n2552));
  andx g2512(.a(n679), .b(n431), .O(n2553));
  andx g2513(.a(n2553), .b(n2552), .O(n2554));
  andx g2514(.a(n2554), .b(n2311), .O(n2555));
  andx g2515(.a(n2555), .b(n2551), .O(n2556));
  orx  g2516(.a(n2556), .b(n2549), .O(n2557));
  orx  g2517(.a(n2557), .b(n2543), .O(n2558));
  andx g2518(.a(n1766), .b(n909), .O(n2559));
  andx g2519(.a(n2559), .b(n2482), .O(n2560));
  andx g2520(.a(n2560), .b(n2480), .O(n2561));
  andx g2521(.a(n2561), .b(n730), .O(n2562));
  andx g2522(.a(n1758), .b(n566), .O(n2563));
  andx g2523(.a(n404), .b(n68), .O(n2564));
  andx g2524(.a(n2564), .b(n2563), .O(n2565));
  andx g2525(.a(n2030), .b(n1976), .O(n2566));
  andx g2526(.a(n2566), .b(n869), .O(n2567));
  andx g2527(.a(n2567), .b(n2565), .O(n2568));
  andx g2528(.a(n2568), .b(n2216), .O(n2569));
  orx  g2529(.a(n2569), .b(n2562), .O(n2570));
  andx g2530(.a(n1056), .b(n1695), .O(n2571));
  andx g2531(.a(n2303), .b(n855), .O(n2572));
  andx g2532(.a(n2572), .b(n1786), .O(n2573));
  andx g2533(.a(n2032), .b(n117), .O(n2574));
  andx g2534(.a(n2209), .b(n459), .O(n2575));
  andx g2535(.a(n2575), .b(n2574), .O(n2576));
  andx g2536(.a(n2576), .b(n2573), .O(n2577));
  andx g2537(.a(n2577), .b(n2571), .O(n2578));
  andx g2538(.a(n459), .b(n268), .O(n2579));
  andx g2539(.a(n2579), .b(n2210), .O(n2580));
  andx g2540(.a(n1848), .b(n1333), .O(n2581));
  andx g2541(.a(n2348), .b(n127), .O(n2582));
  andx g2542(.a(n2582), .b(n2581), .O(n2583));
  andx g2543(.a(n2583), .b(n2580), .O(n2584));
  andx g2544(.a(n2584), .b(n1844), .O(n2585));
  orx  g2545(.a(n2585), .b(n2578), .O(n2586));
  orx  g2546(.a(n2586), .b(n2570), .O(n2587));
  orx  g2547(.a(n2587), .b(n2558), .O(n2588));
  andx g2548(.a(n2039), .b(n1766), .O(n2589));
  andx g2549(.a(n2032), .b(n536), .O(n2590));
  andx g2550(.a(n268), .b(n77), .O(n2591));
  andx g2551(.a(n2591), .b(n2259), .O(n2592));
  andx g2552(.a(n2592), .b(n2590), .O(n2593));
  andx g2553(.a(n2593), .b(n2589), .O(n2594));
  andx g2554(.a(n2461), .b(n430), .O(n2595));
  andx g2555(.a(n2595), .b(n2563), .O(n2596));
  andx g2556(.a(n1344), .b(n428), .O(n2597));
  andx g2557(.a(n2597), .b(n577), .O(n2598));
  andx g2558(.a(n2598), .b(n2596), .O(n2599));
  andx g2559(.a(n2599), .b(n730), .O(n2600));
  orx  g2560(.a(n2600), .b(n2594), .O(n2601));
  andx g2561(.a(n2544), .b(n895), .O(n2602));
  andx g2562(.a(n2602), .b(n2461), .O(n2603));
  andx g2563(.a(n171), .b(n57), .O(n2604));
  andx g2564(.a(n1758), .b(n589), .O(n2605));
  andx g2565(.a(n2605), .b(n2604), .O(n2606));
  andx g2566(.a(n2606), .b(n2603), .O(n2607));
  andx g2567(.a(n2607), .b(n1651), .O(n2608));
  andx g2568(.a(n136), .b(n277), .O(n2609));
  andx g2569(.a(n268), .b(n171), .O(n2610));
  andx g2570(.a(n2610), .b(n2380), .O(n2611));
  andx g2571(.a(n2611), .b(n2609), .O(n2612));
  andx g2572(.a(n2612), .b(n2551), .O(n2613));
  orx  g2573(.a(n2613), .b(n2608), .O(n2614));
  orx  g2574(.a(n2614), .b(n2601), .O(n2615));
  andx g2575(.a(n2045), .b(n93), .O(n2616));
  andx g2576(.a(n1921), .b(n273), .O(n2617));
  andx g2577(.a(n2617), .b(n932), .O(n2618));
  andx g2578(.a(n2618), .b(n2616), .O(n2619));
  andx g2579(.a(n2619), .b(n2453), .O(n2620));
  andx g2580(.a(n1044), .b(n88), .O(n2621));
  andx g2581(.a(n428), .b(n64), .O(n2622));
  andx g2582(.a(n1758), .b(n53), .O(n2623));
  andx g2583(.a(n2623), .b(n2481), .O(n2624));
  andx g2584(.a(n2624), .b(n2622), .O(n2625));
  andx g2585(.a(n2625), .b(n2621), .O(n2626));
  orx  g2586(.a(n2626), .b(n2620), .O(n2627));
  andx g2587(.a(n1844), .b(n268), .O(n2628));
  andx g2588(.a(n214), .b(n59), .O(n2629));
  andx g2589(.a(n1921), .b(n1344), .O(n2630));
  andx g2590(.a(n2630), .b(n2629), .O(n2631));
  andx g2591(.a(n277), .b(n212), .O(n2632));
  andx g2592(.a(n2632), .b(n536), .O(n2633));
  andx g2593(.a(n2633), .b(n205), .O(n2634));
  andx g2594(.a(n2634), .b(n2631), .O(n2635));
  andx g2595(.a(n2635), .b(n2628), .O(n2636));
  andx g2596(.a(n2461), .b(n164), .O(n2637));
  andx g2597(.a(n1758), .b(n545), .O(n2638));
  andx g2598(.a(n2638), .b(n2637), .O(n2639));
  andx g2599(.a(n935), .b(n60), .O(n2640));
  andx g2600(.a(n1951), .b(n2640), .O(n2641));
  andx g2601(.a(n2641), .b(n2639), .O(n2642));
  andx g2602(.a(n2642), .b(n923), .O(n2643));
  orx  g2603(.a(n2643), .b(n2636), .O(n2644));
  orx  g2604(.a(n2644), .b(n2627), .O(n2645));
  orx  g2605(.a(n2645), .b(n2615), .O(n2646));
  orx  g2606(.a(n2646), .b(n2588), .O(n2647));
  orx  g2607(.a(n2647), .b(n2528), .O(n2648));
  andx g2608(.a(n566), .b(n273), .O(n2649));
  andx g2609(.a(n2649), .b(n856), .O(n2650));
  andx g2610(.a(n1694), .b(n1344), .O(n2651));
  andx g2611(.a(n2651), .b(n2015), .O(n2652));
  andx g2612(.a(n2652), .b(n2650), .O(n2653));
  andx g2613(.a(n2653), .b(n2039), .O(n2654));
  andx g2614(.a(n1844), .b(n1811), .O(n2655));
  andx g2615(.a(n2016), .b(n136), .O(n2656));
  andx g2616(.a(n2300), .b(n72), .O(n2657));
  andx g2617(.a(n2303), .b(n2258), .O(n2658));
  andx g2618(.a(n2658), .b(n2657), .O(n2659));
  andx g2619(.a(n2659), .b(n2656), .O(n2660));
  andx g2620(.a(n2660), .b(n2655), .O(n2661));
  orx  g2621(.a(n2661), .b(n2654), .O(n2662));
  andx g2622(.a(n2348), .b(n2231), .O(n2663));
  andx g2623(.a(n2663), .b(n895), .O(n2664));
  andx g2624(.a(n254), .b(n58), .O(n2665));
  andx g2625(.a(n2665), .b(n460), .O(n2666));
  andx g2626(.a(n2666), .b(n2664), .O(n2667));
  andx g2627(.a(n2667), .b(n923), .O(n2668));
  andx g2628(.a(n2032), .b(n61), .O(n2669));
  andx g2629(.a(n1811), .b(n428), .O(n2670));
  andx g2630(.a(n268), .b(n120), .O(n2671));
  andx g2631(.a(n2671), .b(n2670), .O(n2672));
  andx g2632(.a(n2672), .b(n2669), .O(n2673));
  andx g2633(.a(n2673), .b(n2011), .O(n2674));
  orx  g2634(.a(n2674), .b(n2668), .O(n2675));
  orx  g2635(.a(n2675), .b(n2662), .O(n2676));
  andx g2636(.a(n1780), .b(n206), .O(n2677));
  andx g2637(.a(n2677), .b(n2520), .O(n2678));
  andx g2638(.a(n2678), .b(n2604), .O(n2679));
  andx g2639(.a(n2679), .b(n2435), .O(n2680));
  orx  g2640(.a(n2680), .b(n1574), .O(n2681));
  andx g2641(.a(n42), .b(n52), .O(n2682));
  andx g2642(.a(n2682), .b(n381), .O(n2683));
  andx g2643(.a(n2683), .b(n677), .O(n2684));
  andx g2644(.a(n2243), .b(n1667), .O(n2685));
  andx g2645(.a(n2685), .b(n1666), .O(n2686));
  andx g2646(.a(n2686), .b(n2684), .O(n2687));
  andx g2647(.a(n1758), .b(n206), .O(n2688));
  andx g2648(.a(n2688), .b(n2637), .O(n2689));
  andx g2649(.a(n58), .b(n214), .O(n2690));
  andx g2650(.a(n2538), .b(n119), .O(n2691));
  andx g2651(.a(n2691), .b(n2690), .O(n2692));
  andx g2652(.a(n2692), .b(n2689), .O(n2693));
  andx g2653(.a(n2693), .b(n677), .O(n2694));
  orx  g2654(.a(n2694), .b(n2687), .O(n2695));
  orx  g2655(.a(n2695), .b(n2681), .O(n2696));
  andx g2656(.a(n922), .b(n127), .O(n2697));
  andx g2657(.a(n2231), .b(n1694), .O(n2698));
  andx g2658(.a(n2698), .b(n895), .O(n2699));
  andx g2659(.a(n2030), .b(n171), .O(n2700));
  andx g2660(.a(n566), .b(n65), .O(n2701));
  andx g2661(.a(n2701), .b(n2700), .O(n2702));
  andx g2662(.a(n2702), .b(n2699), .O(n2703));
  andx g2663(.a(n2703), .b(n2697), .O(n2704));
  andx g2664(.a(n93), .b(n277), .O(n2705));
  andx g2665(.a(n2705), .b(n117), .O(n2706));
  andx g2666(.a(n1758), .b(n369), .O(n2707));
  andx g2667(.a(n171), .b(n120), .O(n2708));
  andx g2668(.a(n2708), .b(n2707), .O(n2709));
  andx g2669(.a(n2709), .b(n2706), .O(n2710));
  andx g2670(.a(n2710), .b(n2028), .O(n2711));
  orx  g2671(.a(n2711), .b(n2704), .O(n2712));
  andx g2672(.a(n229), .b(pi07), .O(n2713));
  andx g2673(.a(n2231), .b(n1766), .O(n2714));
  andx g2674(.a(n345), .b(n68), .O(n2715));
  andx g2675(.a(n2715), .b(n2714), .O(n2716));
  andx g2676(.a(n2716), .b(n2713), .O(n2717));
  andx g2677(.a(n2717), .b(n1609), .O(n2718));
  andx g2678(.a(n2689), .b(n2311), .O(n2719));
  andx g2679(.a(n2719), .b(n2621), .O(n2720));
  orx  g2680(.a(n2720), .b(n2718), .O(n2721));
  orx  g2681(.a(n2721), .b(n2712), .O(n2722));
  orx  g2682(.a(n2722), .b(n2696), .O(n2723));
  orx  g2683(.a(n2723), .b(n2676), .O(n2724));
  andx g2684(.a(n1321), .b(n1695), .O(n2725));
  andx g2685(.a(n2401), .b(n2258), .O(n2726));
  andx g2686(.a(n277), .b(n91), .O(n2727));
  andx g2687(.a(n2727), .b(n1832), .O(n2728));
  andx g2688(.a(n2728), .b(n1758), .O(n2729));
  andx g2689(.a(n2729), .b(n2726), .O(n2730));
  andx g2690(.a(n2730), .b(n2725), .O(n2731));
  andx g2691(.a(n909), .b(n164), .O(n2732));
  andx g2692(.a(n1811), .b(n545), .O(n2733));
  andx g2693(.a(n2733), .b(n2732), .O(n2734));
  andx g2694(.a(n2734), .b(n286), .O(n2735));
  andx g2695(.a(n2735), .b(n1652), .O(n2736));
  orx  g2696(.a(n2736), .b(n2731), .O(n2737));
  andx g2697(.a(n2688), .b(n2595), .O(n2738));
  andx g2698(.a(n2738), .b(n2692), .O(n2739));
  andx g2699(.a(n2739), .b(n730), .O(n2740));
  andx g2700(.a(n2231), .b(n1243), .O(n2741));
  andx g2701(.a(n345), .b(n182), .O(n2742));
  andx g2702(.a(n2742), .b(n1786), .O(n2743));
  andx g2703(.a(n2743), .b(n105), .O(n2744));
  andx g2704(.a(n2744), .b(n2741), .O(n2745));
  orx  g2705(.a(n2745), .b(n2740), .O(n2746));
  orx  g2706(.a(n2746), .b(n2737), .O(n2747));
  andx g2707(.a(n1148), .b(n397), .O(n2748));
  andx g2708(.a(n2748), .b(n1833), .O(n2749));
  andx g2709(.a(n2749), .b(n1795), .O(n2750));
  andx g2710(.a(n2750), .b(n2279), .O(n2751));
  andx g2711(.a(n1766), .b(n228), .O(n2752));
  andx g2712(.a(n2752), .b(n433), .O(n2753));
  andx g2713(.a(n2753), .b(n1850), .O(n2754));
  andx g2714(.a(n2754), .b(n2039), .O(n2755));
  orx  g2715(.a(n2755), .b(n2751), .O(n2756));
  andx g2716(.a(n943), .b(n41), .O(n2757));
  andx g2717(.a(n668), .b(n2698), .O(n2758));
  andx g2718(.a(n2758), .b(n495), .O(n2759));
  andx g2719(.a(n2759), .b(n2757), .O(n2760));
  andx g2720(.a(n2303), .b(n204), .O(n2761));
  andx g2721(.a(n2761), .b(n1766), .O(n2762));
  andx g2722(.a(n1344), .b(n57), .O(n2763));
  andx g2723(.a(n1999), .b(n364), .O(n2764));
  andx g2724(.a(n2764), .b(n2763), .O(n2765));
  andx g2725(.a(n2765), .b(n2762), .O(n2766));
  andx g2726(.a(n2766), .b(n2427), .O(n2767));
  orx  g2727(.a(n2767), .b(n2760), .O(n2768));
  orx  g2728(.a(n2768), .b(n2756), .O(n2769));
  orx  g2729(.a(n2769), .b(n2747), .O(n2770));
  andx g2730(.a(n2738), .b(n2311), .O(n2771));
  andx g2731(.a(n2771), .b(n1565), .O(n2772));
  andx g2732(.a(n1243), .b(n41), .O(n2773));
  andx g2733(.a(n589), .b(n381), .O(n2774));
  andx g2734(.a(n2461), .b(n238), .O(n2775));
  andx g2735(.a(n2775), .b(n2774), .O(n2776));
  andx g2736(.a(n2776), .b(n1059), .O(n2777));
  andx g2737(.a(n2777), .b(n2773), .O(n2778));
  orx  g2738(.a(n2778), .b(n2772), .O(n2779));
  andx g2739(.a(n2461), .b(n119), .O(n2780));
  andx g2740(.a(n2780), .b(n2563), .O(n2781));
  andx g2741(.a(n802), .b(n108), .O(n2782));
  andx g2742(.a(n2782), .b(n2781), .O(n2783));
  andx g2743(.a(n2783), .b(n943), .O(n2784));
  andx g2744(.a(n59), .b(n1687), .O(n2785));
  andx g2745(.a(n2785), .b(n1198), .O(n2786));
  andx g2746(.a(n1780), .b(n1759), .O(n2787));
  andx g2747(.a(n2787), .b(n2786), .O(n2788));
  andx g2748(.a(n2788), .b(n1700), .O(n2789));
  andx g2749(.a(n2789), .b(n1195), .O(n2790));
  orx  g2750(.a(n2790), .b(n2784), .O(n2791));
  orx  g2751(.a(n2791), .b(n2779), .O(n2792));
  andx g2752(.a(n323), .b(n68), .O(n2793));
  andx g2753(.a(n2793), .b(n2649), .O(n2794));
  andx g2754(.a(n2794), .b(n2652), .O(n2795));
  andx g2755(.a(n2795), .b(n1844), .O(n2796));
  andx g2756(.a(n364), .b(n72), .O(n2797));
  andx g2757(.a(n2797), .b(n1080), .O(n2798));
  andx g2758(.a(n2798), .b(n2495), .O(n2799));
  andx g2759(.a(n2799), .b(n2655), .O(n2800));
  orx  g2760(.a(n2800), .b(n2796), .O(n2801));
  andx g2761(.a(n2550), .b(n979), .O(n2802));
  andx g2762(.a(n2045), .b(n56), .O(n2803));
  andx g2763(.a(n1832), .b(n1344), .O(n2804));
  andx g2764(.a(n2804), .b(n2803), .O(n2805));
  andx g2765(.a(n2805), .b(n2802), .O(n2806));
  andx g2766(.a(n2806), .b(n2039), .O(n2807));
  andx g2767(.a(n1831), .b(n895), .O(n2808));
  andx g2768(.a(n2808), .b(n2231), .O(n2809));
  andx g2769(.a(n2804), .b(n1604), .O(n2810));
  andx g2770(.a(n2810), .b(n2809), .O(n2811));
  andx g2771(.a(n2811), .b(n2697), .O(n2812));
  orx  g2772(.a(n2812), .b(n2807), .O(n2813));
  orx  g2773(.a(n2813), .b(n2801), .O(n2814));
  orx  g2774(.a(n2814), .b(n2792), .O(n2815));
  orx  g2775(.a(n2815), .b(n2770), .O(n2816));
  orx  g2776(.a(n2816), .b(n2724), .O(n2817));
  orx  g2777(.a(n2817), .b(n2648), .O(n2818));
  andx g2778(.a(n2016), .b(n1610), .O(n2819));
  andx g2779(.a(n1838), .b(n431), .O(n2820));
  andx g2780(.a(n2820), .b(n2819), .O(n2821));
  andx g2781(.a(n2821), .b(n2281), .O(n2822));
  andx g2782(.a(n2822), .b(n2309), .O(n2823));
  andx g2783(.a(n943), .b(pi07), .O(n2824));
  andx g2784(.a(n42), .b(n41), .O(n2825));
  andx g2785(.a(n2825), .b(n323), .O(n2826));
  andx g2786(.a(n1832), .b(n1688), .O(n2827));
  andx g2787(.a(n2827), .b(n2826), .O(n2828));
  andx g2788(.a(n2828), .b(n2402), .O(n2829));
  andx g2789(.a(n2829), .b(n2824), .O(n2830));
  orx  g2790(.a(n2830), .b(n2823), .O(n2831));
  andx g2791(.a(n41), .b(n1687), .O(n2832));
  andx g2792(.a(n2832), .b(n1706), .O(n2833));
  andx g2793(.a(n2833), .b(n494), .O(n2834));
  andx g2794(.a(n2637), .b(n1544), .O(n2835));
  andx g2795(.a(n2835), .b(n2834), .O(n2836));
  andx g2796(.a(n2836), .b(n1044), .O(n2837));
  andx g2797(.a(n1942), .b(n1831), .O(n2838));
  andx g2798(.a(n2838), .b(n2461), .O(n2839));
  andx g2799(.a(n2135), .b(n494), .O(n2840));
  andx g2800(.a(n2840), .b(n1544), .O(n2841));
  andx g2801(.a(n2841), .b(n2839), .O(n2842));
  andx g2802(.a(n2842), .b(n677), .O(n2843));
  orx  g2803(.a(n2843), .b(n2837), .O(n2844));
  orx  g2804(.a(n2844), .b(n2831), .O(n2845));
  andx g2805(.a(n668), .b(n248), .O(n2846));
  andx g2806(.a(n2846), .b(n196), .O(n2847));
  andx g2807(.a(n932), .b(n1000), .O(n2848));
  orx  g2808(.a(n2848), .b(n2847), .O(n2849));
  andx g2809(.a(n228), .b(n63), .O(n2850));
  andx g2810(.a(n2850), .b(n125), .O(n2851));
  andx g2811(.a(n2851), .b(n2264), .O(n2852));
  andx g2812(.a(n2474), .b(n450), .O(n2853));
  orx  g2813(.a(n2853), .b(n2852), .O(n2854));
  orx  g2814(.a(n2854), .b(n2849), .O(n2855));
  orx  g2815(.a(n2855), .b(n2845), .O(n2856));
  andx g2816(.a(n92), .b(n249), .O(n2857));
  andx g2817(.a(n2857), .b(n1075), .O(n2858));
  andx g2818(.a(n2135), .b(n1786), .O(n2859));
  andx g2819(.a(n2859), .b(n2858), .O(n2860));
  andx g2820(.a(n2832), .b(n2595), .O(n2861));
  andx g2821(.a(n494), .b(n431), .O(n2862));
  andx g2822(.a(n2862), .b(n1544), .O(n2863));
  andx g2823(.a(n2863), .b(n2861), .O(n2864));
  andx g2824(.a(n2864), .b(n1564), .O(n2865));
  orx  g2825(.a(n2865), .b(n2860), .O(n2866));
  andx g2826(.a(n1811), .b(n1344), .O(n2867));
  andx g2827(.a(n718), .b(n72), .O(n2868));
  andx g2828(.a(n2868), .b(n2867), .O(n2869));
  andx g2829(.a(n2256), .b(n1976), .O(n2870));
  andx g2830(.a(n2870), .b(n1220), .O(n2871));
  andx g2831(.a(n2871), .b(n2869), .O(n2872));
  andx g2832(.a(n2872), .b(n2039), .O(n2873));
  andx g2833(.a(n2673), .b(n2040), .O(n2874));
  orx  g2834(.a(n2874), .b(n2873), .O(n2875));
  orx  g2835(.a(n2875), .b(n2866), .O(n2876));
  andx g2836(.a(n2333), .b(n1831), .O(n2877));
  andx g2837(.a(n2231), .b(n323), .O(n2878));
  andx g2838(.a(n2401), .b(n1832), .O(n2879));
  andx g2839(.a(n2879), .b(n2878), .O(n2880));
  andx g2840(.a(n2880), .b(n2877), .O(n2881));
  andx g2841(.a(n2881), .b(n2824), .O(n2882));
  andx g2842(.a(n2231), .b(n1786), .O(n2883));
  andx g2843(.a(n2883), .b(n430), .O(n2884));
  andx g2844(.a(n2884), .b(n2863), .O(n2885));
  andx g2845(.a(n2885), .b(n1628), .O(n2886));
  orx  g2846(.a(n2886), .b(n2882), .O(n2887));
  andx g2847(.a(n2012), .b(n545), .O(n2888));
  andx g2848(.a(n2888), .b(n164), .O(n2889));
  andx g2849(.a(n2231), .b(n1780), .O(n2890));
  andx g2850(.a(n2890), .b(n2604), .O(n2891));
  andx g2851(.a(n2891), .b(n2889), .O(n2892));
  andx g2852(.a(n2892), .b(n2697), .O(n2893));
  andx g2853(.a(n1773), .b(n228), .O(n2894));
  andx g2854(.a(n2894), .b(n895), .O(n2895));
  andx g2855(.a(n1344), .b(n56), .O(n2896));
  andx g2856(.a(n1999), .b(n1694), .O(n2897));
  andx g2857(.a(n2897), .b(n2896), .O(n2898));
  andx g2858(.a(n2898), .b(n2895), .O(n2899));
  andx g2859(.a(n2899), .b(n2571), .O(n2900));
  orx  g2860(.a(n2900), .b(n2893), .O(n2901));
  orx  g2861(.a(n2901), .b(n2887), .O(n2902));
  orx  g2862(.a(n2902), .b(n2876), .O(n2903));
  orx  g2863(.a(n2903), .b(n2856), .O(n2904));
  andx g2864(.a(n2461), .b(n1758), .O(n2905));
  andx g2865(.a(n2905), .b(n1831), .O(n2906));
  andx g2866(.a(n2906), .b(n2598), .O(n2907));
  andx g2867(.a(n2907), .b(n2232), .O(n2908));
  andx g2868(.a(n1688), .b(n566), .O(n2909));
  andx g2869(.a(n2461), .b(n53), .O(n2910));
  andx g2870(.a(n2910), .b(n2909), .O(n2911));
  andx g2871(.a(n406), .b(n108), .O(n2912));
  andx g2872(.a(n2912), .b(n2911), .O(n2913));
  andx g2873(.a(n2913), .b(n943), .O(n2914));
  orx  g2874(.a(n2914), .b(n2908), .O(n2915));
  andx g2875(.a(n2357), .b(n2258), .O(n2916));
  andx g2876(.a(n536), .b(n278), .O(n2917));
  andx g2877(.a(n369), .b(n264), .O(n2918));
  andx g2878(.a(n2918), .b(n2917), .O(n2919));
  andx g2879(.a(n2919), .b(n2916), .O(n2920));
  andx g2880(.a(n2920), .b(n2655), .O(n2921));
  andx g2881(.a(n65), .b(n75), .O(n2922));
  andx g2882(.a(n2733), .b(n1198), .O(n2923));
  andx g2883(.a(n2923), .b(n2922), .O(n2924));
  andx g2884(.a(n2924), .b(n778), .O(n2925));
  orx  g2885(.a(n2925), .b(n2921), .O(n2926));
  orx  g2886(.a(n2926), .b(n2915), .O(n2927));
  andx g2887(.a(n2231), .b(n566), .O(n2928));
  andx g2888(.a(n2928), .b(n545), .O(n2929));
  andx g2889(.a(n2251), .b(n1108), .O(n2930));
  andx g2890(.a(n2930), .b(n2929), .O(n2931));
  andx g2891(.a(n2931), .b(n2697), .O(n2932));
  andx g2892(.a(n566), .b(n459), .O(n2933));
  andx g2893(.a(n2933), .b(n273), .O(n2934));
  andx g2894(.a(n2032), .b(n136), .O(n2935));
  andx g2895(.a(n127), .b(n104), .O(n2936));
  andx g2896(.a(n2936), .b(n2935), .O(n2937));
  andx g2897(.a(n2937), .b(n2934), .O(n2938));
  andx g2898(.a(n2938), .b(n2028), .O(n2939));
  orx  g2899(.a(n2939), .b(n2932), .O(n2940));
  andx g2900(.a(n2461), .b(n1688), .O(n2941));
  andx g2901(.a(n2941), .b(n895), .O(n2942));
  andx g2902(.a(n2862), .b(n2490), .O(n2943));
  andx g2903(.a(n2943), .b(n2942), .O(n2944));
  andx g2904(.a(n2944), .b(n975), .O(n2945));
  andx g2905(.a(n1610), .b(n329), .O(n2946));
  andx g2906(.a(n1786), .b(n566), .O(n2947));
  andx g2907(.a(n2947), .b(n2946), .O(n2948));
  andx g2908(.a(n2209), .b(n65), .O(n2949));
  andx g2909(.a(n2949), .b(n1544), .O(n2950));
  andx g2910(.a(n2950), .b(n2948), .O(n2951));
  andx g2911(.a(n2951), .b(n975), .O(n2952));
  orx  g2912(.a(n2952), .b(n2945), .O(n2953));
  orx  g2913(.a(n2953), .b(n2940), .O(n2954));
  orx  g2914(.a(n2954), .b(n2927), .O(n2955));
  andx g2915(.a(n437), .b(pi29), .O(n2956));
  andx g2916(.a(n2956), .b(n584), .O(n2957));
  andx g2917(.a(n2957), .b(n196), .O(n2958));
  andx g2918(.a(n1768), .b(n2665), .O(n2959));
  andx g2919(.a(n545), .b(n397), .O(n2960));
  andx g2920(.a(n2960), .b(n2115), .O(n2961));
  andx g2921(.a(n2961), .b(n2959), .O(n2962));
  orx  g2922(.a(n2962), .b(n2958), .O(n2963));
  andx g2923(.a(pi07), .b(n1687), .O(n2964));
  andx g2924(.a(n2964), .b(n1786), .O(n2965));
  andx g2925(.a(n2965), .b(n2858), .O(n2966));
  andx g2926(.a(n396), .b(n80), .O(n2967));
  andx g2927(.a(n1832), .b(n199), .O(n2968));
  andx g2928(.a(n2968), .b(n756), .O(n2969));
  andx g2929(.a(n2969), .b(n2967), .O(n2970));
  orx  g2930(.a(n2970), .b(n2966), .O(n2971));
  orx  g2931(.a(n2971), .b(n2963), .O(n2972));
  andx g2932(.a(n2012), .b(n397), .O(n2973));
  andx g2933(.a(n2973), .b(n895), .O(n2974));
  andx g2934(.a(pi29), .b(n56), .O(n2975));
  andx g2935(.a(n2975), .b(n2032), .O(n2976));
  andx g2936(.a(n2030), .b(n1832), .O(n2977));
  andx g2937(.a(n2977), .b(n2976), .O(n2978));
  andx g2938(.a(n2978), .b(n2974), .O(n2979));
  andx g2939(.a(n2979), .b(n2215), .O(n2980));
  andx g2940(.a(n2231), .b(n1838), .O(n2981));
  andx g2941(.a(n2981), .b(n545), .O(n2982));
  andx g2942(.a(n213), .b(n104), .O(n2983));
  andx g2943(.a(n2401), .b(n68), .O(n2984));
  andx g2944(.a(n2984), .b(n2983), .O(n2985));
  andx g2945(.a(n2985), .b(n2982), .O(n2986));
  andx g2946(.a(n2986), .b(n923), .O(n2987));
  orx  g2947(.a(n2987), .b(n2980), .O(n2988));
  andx g2948(.a(n2428), .b(n254), .O(n2989));
  andx g2949(.a(n2184), .b(n1780), .O(n2990));
  andx g2950(.a(n2990), .b(n2989), .O(n2991));
  andx g2951(.a(n2991), .b(n908), .O(n2992));
  andx g2952(.a(n1688), .b(n1503), .O(n2993));
  andx g2953(.a(n2993), .b(n1766), .O(n2994));
  andx g2954(.a(n2994), .b(n286), .O(n2995));
  andx g2955(.a(n2995), .b(n778), .O(n2996));
  orx  g2956(.a(n2996), .b(n2992), .O(n2997));
  orx  g2957(.a(n2997), .b(n2988), .O(n2998));
  orx  g2958(.a(n2998), .b(n2972), .O(n2999));
  orx  g2959(.a(n2999), .b(n2955), .O(n3000));
  orx  g2960(.a(n3000), .b(n2904), .O(n3001));
  andx g2961(.a(n895), .b(n153), .O(n3002));
  andx g2962(.a(n3002), .b(n2488), .O(n3003));
  andx g2963(.a(n735), .b(n589), .O(n3004));
  andx g2964(.a(n3004), .b(n2311), .O(n3005));
  andx g2965(.a(n3005), .b(n3003), .O(n3006));
  andx g2966(.a(n3006), .b(n975), .O(n3007));
  andx g2967(.a(n329), .b(n119), .O(n3008));
  andx g2968(.a(n1766), .b(n1758), .O(n3009));
  andx g2969(.a(n3009), .b(n3008), .O(n3010));
  andx g2970(.a(n2538), .b(n589), .O(n3011));
  andx g2971(.a(n3011), .b(n2690), .O(n3012));
  andx g2972(.a(n3012), .b(n3010), .O(n3013));
  andx g2973(.a(n3013), .b(n730), .O(n3014));
  orx  g2974(.a(n3014), .b(n3007), .O(n3015));
  andx g2975(.a(n943), .b(n52), .O(n3016));
  andx g2976(.a(n909), .b(n573), .O(n3017));
  andx g2977(.a(n902), .b(n428), .O(n3018));
  andx g2978(.a(n41), .b(pi37), .O(n3019));
  andx g2979(.a(n3019), .b(n1758), .O(n3020));
  andx g2980(.a(n3020), .b(n3018), .O(n3021));
  andx g2981(.a(n3021), .b(n3017), .O(n3022));
  andx g2982(.a(n3022), .b(n3016), .O(n3023));
  andx g2983(.a(n1831), .b(n53), .O(n3024));
  andx g2984(.a(n3024), .b(n2231), .O(n3025));
  andx g2985(.a(n1786), .b(n76), .O(n3026));
  andx g2986(.a(n3026), .b(n588), .O(n3027));
  andx g2987(.a(n3027), .b(n3025), .O(n3028));
  andx g2988(.a(n3028), .b(n677), .O(n3029));
  orx  g2989(.a(n3029), .b(n3023), .O(n3030));
  orx  g2990(.a(n3030), .b(n3015), .O(n3031));
  andx g2991(.a(n182), .b(n89), .O(n3032));
  andx g2992(.a(n3032), .b(n2595), .O(n3033));
  andx g2993(.a(n3033), .b(n105), .O(n3034));
  andx g2994(.a(n3034), .b(n1348), .O(n3035));
  andx g2995(.a(n171), .b(n60), .O(n3036));
  andx g2996(.a(n2461), .b(n307), .O(n3037));
  andx g2997(.a(n3037), .b(n2605), .O(n3038));
  andx g2998(.a(n3038), .b(n3036), .O(n3039));
  andx g2999(.a(n3039), .b(n2459), .O(n3040));
  orx  g3000(.a(n3040), .b(n3035), .O(n3041));
  andx g3001(.a(n1976), .b(n369), .O(n3042));
  andx g3002(.a(n3042), .b(n2340), .O(n3043));
  andx g3003(.a(n3043), .b(n2916), .O(n3044));
  andx g3004(.a(n3044), .b(n2494), .O(n3045));
  andx g3005(.a(n2209), .b(n1344), .O(n3046));
  andx g3006(.a(n3046), .b(n61), .O(n3047));
  andx g3007(.a(n1848), .b(n68), .O(n3048));
  andx g3008(.a(n3048), .b(n2582), .O(n3049));
  andx g3009(.a(n3049), .b(n3047), .O(n3050));
  andx g3010(.a(n3050), .b(n2628), .O(n3051));
  orx  g3011(.a(n3051), .b(n3045), .O(n3052));
  orx  g3012(.a(n3052), .b(n3041), .O(n3053));
  orx  g3013(.a(n3053), .b(n3031), .O(n3054));
  andx g3014(.a(n41), .b(n52), .O(n3055));
  andx g3015(.a(n3055), .b(n381), .O(n3056));
  andx g3016(.a(n3056), .b(n2461), .O(n3057));
  andx g3017(.a(n2949), .b(n163), .O(n3058));
  andx g3018(.a(n3058), .b(n3057), .O(n3059));
  andx g3019(.a(n3059), .b(n1044), .O(n3060));
  andx g3020(.a(n2589), .b(n2306), .O(n3061));
  orx  g3021(.a(n3061), .b(n3060), .O(n3062));
  andx g3022(.a(n204), .b(n58), .O(n3063));
  andx g3023(.a(n2461), .b(n199), .O(n3064));
  andx g3024(.a(n3064), .b(n3063), .O(n3065));
  andx g3025(.a(n3065), .b(n2877), .O(n3066));
  andx g3026(.a(n3066), .b(n3016), .O(n3067));
  andx g3027(.a(n1786), .b(n545), .O(n3068));
  andx g3028(.a(n3068), .b(n2231), .O(n3069));
  andx g3029(.a(n494), .b(n65), .O(n3070));
  andx g3030(.a(n3070), .b(n1544), .O(n3071));
  andx g3031(.a(n3071), .b(n3069), .O(n3072));
  andx g3032(.a(n3072), .b(n1628), .O(n3073));
  orx  g3033(.a(n3073), .b(n3067), .O(n3074));
  orx  g3034(.a(n3074), .b(n3062), .O(n3075));
  andx g3035(.a(n2727), .b(n171), .O(n3076));
  andx g3036(.a(n120), .b(n104), .O(n3077));
  andx g3037(.a(n3077), .b(n1811), .O(n3078));
  andx g3038(.a(n3078), .b(n3076), .O(n3079));
  andx g3039(.a(n3079), .b(n2725), .O(n3080));
  andx g3040(.a(n1786), .b(n345), .O(n3081));
  andx g3041(.a(n3081), .b(n53), .O(n3082));
  andx g3042(.a(n3082), .b(n105), .O(n3083));
  andx g3043(.a(n3083), .b(n2741), .O(n3084));
  orx  g3044(.a(n3084), .b(n3080), .O(n3085));
  andx g3045(.a(n1148), .b(n273), .O(n3086));
  andx g3046(.a(n1786), .b(n735), .O(n3087));
  andx g3047(.a(n3087), .b(n3086), .O(n3088));
  andx g3048(.a(n2045), .b(n87), .O(n3089));
  andx g3049(.a(n733), .b(n171), .O(n3090));
  andx g3050(.a(n3090), .b(n3089), .O(n3091));
  andx g3051(.a(n3091), .b(n3088), .O(n3092));
  andx g3052(.a(n3092), .b(n2215), .O(n3093));
  andx g3053(.a(n2219), .b(n264), .O(n3094));
  andx g3054(.a(n3094), .b(n2579), .O(n3095));
  andx g3055(.a(n2348), .b(n840), .O(n3096));
  andx g3056(.a(n2300), .b(n1204), .O(n3097));
  andx g3057(.a(n3097), .b(n3096), .O(n3098));
  andx g3058(.a(n3098), .b(n3095), .O(n3099));
  andx g3059(.a(n3099), .b(n2215), .O(n3100));
  orx  g3060(.a(n3100), .b(n3093), .O(n3101));
  orx  g3061(.a(n3101), .b(n3085), .O(n3102));
  orx  g3062(.a(n3102), .b(n3075), .O(n3103));
  orx  g3063(.a(n3103), .b(n3054), .O(n3104));
  andx g3064(.a(n494), .b(n73), .O(n3105));
  andx g3065(.a(n3105), .b(n2890), .O(n3106));
  andx g3066(.a(n3106), .b(n1544), .O(n3107));
  andx g3067(.a(n3107), .b(n2757), .O(n3108));
  andx g3068(.a(n2219), .b(n1838), .O(n3109));
  andx g3069(.a(n3109), .b(n406), .O(n3110));
  andx g3070(.a(n3110), .b(n1211), .O(n3111));
  andx g3071(.a(n3111), .b(n2684), .O(n3112));
  orx  g3072(.a(n3112), .b(n3108), .O(n3113));
  andx g3073(.a(n2516), .b(n1815), .O(n3114));
  andx g3074(.a(n3114), .b(n1343), .O(n3115));
  andx g3075(.a(n3115), .b(n196), .O(n3116));
  andx g3076(.a(n1758), .b(n329), .O(n3117));
  andx g3077(.a(n3117), .b(n1989), .O(n3118));
  andx g3078(.a(n3118), .b(n2095), .O(n3119));
  andx g3079(.a(n3119), .b(n1652), .O(n3120));
  orx  g3080(.a(n3120), .b(n3116), .O(n3121));
  orx  g3081(.a(n3121), .b(n3113), .O(n3122));
  andx g3082(.a(n2832), .b(n2559), .O(n3123));
  andx g3083(.a(n2763), .b(n69), .O(n3124));
  andx g3084(.a(n3124), .b(n3123), .O(n3125));
  andx g3085(.a(n3125), .b(n1651), .O(n3126));
  andx g3086(.a(n1831), .b(n1148), .O(n3127));
  andx g3087(.a(n3127), .b(n2461), .O(n3128));
  andx g3088(.a(n397), .b(n206), .O(n3129));
  andx g3089(.a(n3129), .b(n2311), .O(n3130));
  andx g3090(.a(n3130), .b(n3128), .O(n3131));
  andx g3091(.a(n3131), .b(n730), .O(n3132));
  orx  g3092(.a(n3132), .b(n3126), .O(n3133));
  andx g3093(.a(n286), .b(n73), .O(n3134));
  andx g3094(.a(n3134), .b(n1000), .O(n3135));
  orx  g3095(.a(n3135), .b(n1546), .O(n3136));
  orx  g3096(.a(n3136), .b(n3133), .O(n3137));
  orx  g3097(.a(n3137), .b(n3122), .O(n3138));
  andx g3098(.a(n164), .b(n1687), .O(n3139));
  andx g3099(.a(n1780), .b(n1198), .O(n3140));
  andx g3100(.a(n3140), .b(n147), .O(n3141));
  andx g3101(.a(n3141), .b(n3139), .O(n3142));
  andx g3102(.a(n3142), .b(n1892), .O(n3143));
  andx g3103(.a(n909), .b(n449), .O(n3144));
  andx g3104(.a(n3144), .b(n3009), .O(n3145));
  andx g3105(.a(n3145), .b(n978), .O(n3146));
  andx g3106(.a(n3146), .b(n1565), .O(n3147));
  orx  g3107(.a(n3147), .b(n3143), .O(n3148));
  andx g3108(.a(n182), .b(n164), .O(n3149));
  andx g3109(.a(n3149), .b(n2714), .O(n3150));
  andx g3110(.a(n3150), .b(n105), .O(n3151));
  andx g3111(.a(n3151), .b(n2509), .O(n3152));
  andx g3112(.a(n1766), .b(n204), .O(n3153));
  andx g3113(.a(n3153), .b(n1810), .O(n3154));
  andx g3114(.a(n3154), .b(n2959), .O(n3155));
  orx  g3115(.a(n3155), .b(n3152), .O(n3156));
  orx  g3116(.a(n3156), .b(n3148), .O(n3157));
  andx g3117(.a(n668), .b(n148), .O(n3158));
  andx g3118(.a(n171), .b(n73), .O(n3159));
  andx g3119(.a(n3159), .b(n1780), .O(n3160));
  andx g3120(.a(n3160), .b(n2967), .O(n3161));
  orx  g3121(.a(n3161), .b(n3158), .O(n3162));
  andx g3122(.a(n2231), .b(n164), .O(n3163));
  andx g3123(.a(n3163), .b(n2677), .O(n3164));
  andx g3124(.a(n3164), .b(n2604), .O(n3165));
  andx g3125(.a(n3165), .b(n2773), .O(n3166));
  andx g3126(.a(n956), .b(n2905), .O(n3167));
  andx g3127(.a(n840), .b(n538), .O(n3168));
  andx g3128(.a(n3168), .b(n2469), .O(n3169));
  andx g3129(.a(n3169), .b(n3167), .O(n3170));
  andx g3130(.a(n3170), .b(n943), .O(n3171));
  orx  g3131(.a(n3171), .b(n3166), .O(n3172));
  orx  g3132(.a(n3172), .b(n3162), .O(n3173));
  orx  g3133(.a(n3173), .b(n3157), .O(n3174));
  orx  g3134(.a(n3174), .b(n3138), .O(n3175));
  orx  g3135(.a(n3175), .b(n3104), .O(n3176));
  orx  g3136(.a(n3176), .b(n3001), .O(n3177));
  orx  g3137(.a(n3177), .b(n2818), .O(n3178));
  orx  g3138(.a(n3178), .b(n2426), .O(po1));
  andx g3139(.a(n44), .b(pi35), .O(n3180));
  andx g3140(.a(n1687), .b(n91), .O(n3181));
  andx g3141(.a(n3181), .b(n67), .O(n3182));
  andx g3142(.a(n3182), .b(n3180), .O(n3183));
  andx g3143(.a(n75), .b(n333), .O(n3184));
  andx g3144(.a(n3184), .b(n431), .O(n3185));
  andx g3145(.a(n3185), .b(n60), .O(n3186));
  invx g3146(.a(pi14), .O(n3187));
  andx g3147(.a(n3187), .b(pi19), .O(n3188));
  andx g3148(.a(pi20), .b(pi17), .O(n3189));
  andx g3149(.a(n3189), .b(n3188), .O(n3190));
  andx g3150(.a(n3190), .b(n3186), .O(n3191));
  andx g3151(.a(n3191), .b(n3183), .O(n3192));
  invx g3152(.a(pi23), .O(n3193));
  andx g3153(.a(n3193), .b(n75), .O(n3194));
  andx g3154(.a(n3194), .b(n107), .O(n3195));
  andx g3155(.a(n42), .b(n151), .O(n3196));
  andx g3156(.a(n3196), .b(n3195), .O(n3197));
  andx g3157(.a(n3197), .b(n644), .O(n3198));
  andx g3158(.a(n46), .b(n63), .O(n3199));
  andx g3159(.a(n44), .b(n87), .O(n3200));
  andx g3160(.a(n3200), .b(n3199), .O(n3201));
  andx g3161(.a(pi14), .b(pi35), .O(n3202));
  andx g3162(.a(n43), .b(n47), .O(n3203));
  andx g3163(.a(n3203), .b(n3202), .O(n3204));
  andx g3164(.a(n3204), .b(n3201), .O(n3205));
  andx g3165(.a(n3205), .b(n3198), .O(n3206));
  orx  g3166(.a(n3206), .b(n3192), .O(n3207));
  andx g3167(.a(n60), .b(pi15), .O(n3208));
  andx g3168(.a(n3208), .b(n333), .O(n3209));
  andx g3169(.a(n3209), .b(n1344), .O(n3210));
  andx g3170(.a(n3210), .b(n3189), .O(n3211));
  andx g3171(.a(pi19), .b(n63), .O(n3212));
  andx g3172(.a(n3212), .b(n313), .O(n3213));
  andx g3173(.a(pi35), .b(n1687), .O(n3214));
  andx g3174(.a(n3214), .b(n91), .O(n3215));
  andx g3175(.a(n3215), .b(n3213), .O(n3216));
  andx g3176(.a(n3216), .b(n3211), .O(n3217));
  andx g3177(.a(n1687), .b(n249), .O(n3218));
  andx g3178(.a(n88), .b(pi35), .O(n3219));
  andx g3179(.a(n3219), .b(n3218), .O(n3220));
  andx g3180(.a(n43), .b(n303), .O(n3221));
  andx g3181(.a(n3221), .b(n48), .O(n3222));
  andx g3182(.a(n3222), .b(n3220), .O(n3223));
  andx g3183(.a(n3185), .b(n42), .O(n3224));
  andx g3184(.a(n3224), .b(n93), .O(n3225));
  andx g3185(.a(n3225), .b(n3223), .O(n3226));
  orx  g3186(.a(n3226), .b(n3217), .O(n3227));
  orx  g3187(.a(n3227), .b(n3207), .O(n3228));
  andx g3188(.a(n3208), .b(n3184), .O(n3229));
  andx g3189(.a(n3229), .b(pi18), .O(n3230));
  andx g3190(.a(n303), .b(n91), .O(n3231));
  andx g3191(.a(n67), .b(n87), .O(n3232));
  andx g3192(.a(n3232), .b(n3231), .O(n3233));
  andx g3193(.a(pi35), .b(n63), .O(n3234));
  andx g3194(.a(n3234), .b(n3189), .O(n3235));
  andx g3195(.a(n3235), .b(n3218), .O(n3236));
  andx g3196(.a(n3236), .b(n3233), .O(n3237));
  andx g3197(.a(n3237), .b(n3230), .O(n3238));
  andx g3198(.a(n3193), .b(n87), .O(n3239));
  andx g3199(.a(pi16), .b(n75), .O(n3240));
  andx g3200(.a(n42), .b(n64), .O(n3241));
  andx g3201(.a(n3241), .b(n3240), .O(n3242));
  andx g3202(.a(n3242), .b(n3239), .O(n3243));
  andx g3203(.a(n533), .b(n41), .O(n3244));
  andx g3204(.a(n3244), .b(n3243), .O(n3245));
  andx g3205(.a(n46), .b(pi35), .O(n3246));
  andx g3206(.a(n3246), .b(n63), .O(n3247));
  andx g3207(.a(n93), .b(n303), .O(n3248));
  andx g3208(.a(n3248), .b(n3203), .O(n3249));
  andx g3209(.a(n3249), .b(n3247), .O(n3250));
  andx g3210(.a(n3250), .b(n3245), .O(n3251));
  orx  g3211(.a(n3251), .b(n3238), .O(n3252));
  andx g3212(.a(n46), .b(n1687), .O(n3253));
  andx g3213(.a(n3253), .b(pi35), .O(n3254));
  andx g3214(.a(n93), .b(n47), .O(n3255));
  andx g3215(.a(n3255), .b(n45), .O(n3256));
  andx g3216(.a(n3256), .b(n3254), .O(n3257));
  andx g3217(.a(n229), .b(n107), .O(n3258));
  andx g3218(.a(n214), .b(n42), .O(n3259));
  andx g3219(.a(n3259), .b(n3258), .O(n3260));
  andx g3220(.a(n212), .b(n64), .O(n3261));
  andx g3221(.a(n3261), .b(pi07), .O(n3262));
  andx g3222(.a(n3262), .b(n3260), .O(n3263));
  andx g3223(.a(n3263), .b(n3257), .O(n3264));
  andx g3224(.a(pi20), .b(n3187), .O(n3265));
  andx g3225(.a(n3265), .b(pi17), .O(n3266));
  andx g3226(.a(n3239), .b(n3184), .O(n3267));
  andx g3227(.a(n3267), .b(n60), .O(n3268));
  andx g3228(.a(n3268), .b(n3266), .O(n3269));
  andx g3229(.a(pi35), .b(n249), .O(n3270));
  andx g3230(.a(n3270), .b(n63), .O(n3271));
  andx g3231(.a(n67), .b(pi19), .O(n3272));
  andx g3232(.a(n3272), .b(n3231), .O(n3273));
  andx g3233(.a(n3273), .b(n3271), .O(n3274));
  andx g3234(.a(n3274), .b(n3269), .O(n3275));
  orx  g3235(.a(n3275), .b(n3264), .O(n3276));
  orx  g3236(.a(n3276), .b(n3252), .O(n3277));
  orx  g3237(.a(n3277), .b(n3228), .O(n3278));
  andx g3238(.a(n3224), .b(n43), .O(n3279));
  andx g3239(.a(n3270), .b(n895), .O(n3280));
  andx g3240(.a(n1773), .b(n48), .O(n3281));
  andx g3241(.a(n3281), .b(n3280), .O(n3282));
  andx g3242(.a(n3282), .b(n3279), .O(n3283));
  andx g3243(.a(n75), .b(pi15), .O(n3284));
  andx g3244(.a(n60), .b(pi18), .O(n3285));
  andx g3245(.a(n3285), .b(pi16), .O(n3286));
  andx g3246(.a(n3286), .b(n3284), .O(n3287));
  andx g3247(.a(n3287), .b(pi07), .O(n3288));
  andx g3248(.a(n1901), .b(n3193), .O(n3289));
  andx g3249(.a(pi35), .b(n303), .O(n3290));
  andx g3250(.a(n3290), .b(n65), .O(n3291));
  andx g3251(.a(n3291), .b(n3289), .O(n3292));
  andx g3252(.a(n3292), .b(n3288), .O(n3293));
  orx  g3253(.a(n3293), .b(n3283), .O(n3294));
  andx g3254(.a(n3259), .b(n3195), .O(n3295));
  andx g3255(.a(n3295), .b(n43), .O(n3296));
  andx g3256(.a(n303), .b(n87), .O(n3297));
  andx g3257(.a(n3297), .b(n3270), .O(n3298));
  andx g3258(.a(n3261), .b(n3199), .O(n3299));
  andx g3259(.a(n3299), .b(n3255), .O(n3300));
  andx g3260(.a(n3300), .b(n3298), .O(n3301));
  andx g3261(.a(n3301), .b(n3296), .O(n3302));
  andx g3262(.a(n3214), .b(n67), .O(n3303));
  andx g3263(.a(n3303), .b(n3222), .O(n3304));
  andx g3264(.a(n60), .b(pi16), .O(n3305));
  andx g3265(.a(n3305), .b(n42), .O(n3306));
  andx g3266(.a(n3306), .b(n229), .O(n3307));
  andx g3267(.a(n73), .b(n41), .O(n3308));
  andx g3268(.a(n3308), .b(n3188), .O(n3309));
  andx g3269(.a(n3309), .b(n3307), .O(n3310));
  andx g3270(.a(n3310), .b(n3304), .O(n3311));
  orx  g3271(.a(n3311), .b(n3302), .O(n3312));
  orx  g3272(.a(n3312), .b(n3294), .O(n3313));
  andx g3273(.a(pi26), .b(n42), .O(n3314));
  andx g3274(.a(n3314), .b(n3258), .O(n3315));
  andx g3275(.a(n3315), .b(n73), .O(n3316));
  andx g3276(.a(n3316), .b(n3257), .O(n3317));
  andx g3277(.a(n333), .b(pi15), .O(n3318));
  andx g3278(.a(n3318), .b(n3306), .O(n3319));
  andx g3279(.a(n91), .b(n63), .O(n3320));
  andx g3280(.a(n3320), .b(n75), .O(n3321));
  andx g3281(.a(n3272), .b(n3239), .O(n3322));
  andx g3282(.a(n3322), .b(n3290), .O(n3323));
  andx g3283(.a(n3323), .b(n3321), .O(n3324));
  andx g3284(.a(n3324), .b(n3319), .O(n3325));
  orx  g3285(.a(n3325), .b(n3317), .O(n3326));
  andx g3286(.a(n3239), .b(n1768), .O(n3327));
  andx g3287(.a(n3327), .b(n855), .O(n3328));
  andx g3288(.a(pi16), .b(pi19), .O(n3329));
  andx g3289(.a(n3329), .b(pi20), .O(n3330));
  andx g3290(.a(n3330), .b(n3229), .O(n3331));
  andx g3291(.a(n3331), .b(pi35), .O(n3332));
  andx g3292(.a(n3332), .b(n3328), .O(n3333));
  andx g3293(.a(n3224), .b(n41), .O(n3334));
  andx g3294(.a(n3334), .b(n3257), .O(n3335));
  orx  g3295(.a(n3335), .b(n3333), .O(n3336));
  orx  g3296(.a(n3336), .b(n3326), .O(n3337));
  orx  g3297(.a(n3337), .b(n3313), .O(n3338));
  orx  g3298(.a(n3338), .b(n3278), .O(n3339));
  andx g3299(.a(n3320), .b(n303), .O(n3340));
  andx g3300(.a(n3214), .b(n164), .O(n3341));
  andx g3301(.a(n3341), .b(n3340), .O(n3342));
  andx g3302(.a(n3342), .b(n3288), .O(n3343));
  andx g3303(.a(n3267), .b(n42), .O(n3344));
  andx g3304(.a(n3344), .b(n43), .O(n3345));
  andx g3305(.a(n88), .b(n303), .O(n3346));
  andx g3306(.a(n3346), .b(n3234), .O(n3347));
  andx g3307(.a(n1689), .b(n48), .O(n3348));
  andx g3308(.a(n3348), .b(n3347), .O(n3349));
  andx g3309(.a(n3349), .b(n3345), .O(n3350));
  orx  g3310(.a(n3350), .b(n3343), .O(n3351));
  andx g3311(.a(n73), .b(pi14), .O(n3352));
  andx g3312(.a(n3352), .b(n3197), .O(n3353));
  andx g3313(.a(n3203), .b(n3180), .O(n3354));
  andx g3314(.a(n1942), .b(n46), .O(n3355));
  andx g3315(.a(n3355), .b(n3354), .O(n3356));
  andx g3316(.a(n3356), .b(n3353), .O(n3357));
  andx g3317(.a(n3184), .b(n107), .O(n3358));
  andx g3318(.a(n3358), .b(n3314), .O(n3359));
  andx g3319(.a(n943), .b(n3359), .O(n3360));
  andx g3320(.a(n3214), .b(n431), .O(n3361));
  andx g3321(.a(n3361), .b(n3360), .O(n3362));
  orx  g3322(.a(n3362), .b(n3357), .O(n3363));
  orx  g3323(.a(n3363), .b(n3351), .O(n3364));
  andx g3324(.a(n1344), .b(n107), .O(n3365));
  andx g3325(.a(n3365), .b(n3196), .O(n3366));
  andx g3326(.a(n47), .b(n1687), .O(n3367));
  andx g3327(.a(n3367), .b(n3202), .O(n3368));
  andx g3328(.a(n43), .b(n46), .O(n3369));
  andx g3329(.a(n3369), .b(n644), .O(n3370));
  andx g3330(.a(n3370), .b(n3368), .O(n3371));
  andx g3331(.a(n3371), .b(n1335), .O(n3372));
  andx g3332(.a(n3372), .b(n3366), .O(n3373));
  andx g3333(.a(n3270), .b(n855), .O(n3374));
  andx g3334(.a(n67), .b(n212), .O(n3375));
  andx g3335(.a(n3375), .b(n73), .O(n3376));
  andx g3336(.a(n3376), .b(n48), .O(n3377));
  andx g3337(.a(n3377), .b(n3374), .O(n3378));
  andx g3338(.a(n3378), .b(n3296), .O(n3379));
  orx  g3339(.a(n3379), .b(n3373), .O(n3380));
  andx g3340(.a(n3358), .b(n3259), .O(n3381));
  andx g3341(.a(n43), .b(n212), .O(n3382));
  andx g3342(.a(n3382), .b(n48), .O(n3383));
  andx g3343(.a(n3383), .b(n3381), .O(n3384));
  andx g3344(.a(n895), .b(n87), .O(n3385));
  andx g3345(.a(n3270), .b(n1758), .O(n3386));
  andx g3346(.a(n3386), .b(n3385), .O(n3387));
  andx g3347(.a(n3387), .b(n3384), .O(n3388));
  andx g3348(.a(n42), .b(n333), .O(n3389));
  andx g3349(.a(n3194), .b(pi16), .O(n3390));
  andx g3350(.a(n3390), .b(n3389), .O(n3391));
  andx g3351(.a(n3391), .b(n93), .O(n3392));
  andx g3352(.a(n855), .b(n87), .O(n3393));
  andx g3353(.a(n88), .b(n533), .O(n3394));
  andx g3354(.a(n3394), .b(n3246), .O(n3395));
  andx g3355(.a(n3395), .b(n3203), .O(n3396));
  andx g3356(.a(n3396), .b(n3393), .O(n3397));
  andx g3357(.a(n3397), .b(n3392), .O(n3398));
  orx  g3358(.a(n3398), .b(n3388), .O(n3399));
  orx  g3359(.a(n3399), .b(n3380), .O(n3400));
  orx  g3360(.a(n3400), .b(n3364), .O(n3401));
  andx g3361(.a(n1942), .b(n75), .O(n3402));
  andx g3362(.a(n42), .b(n3193), .O(n3403));
  andx g3363(.a(n3403), .b(n3402), .O(n3404));
  andx g3364(.a(n3404), .b(pi07), .O(n3405));
  andx g3365(.a(n46), .b(n303), .O(n3406));
  andx g3366(.a(n3406), .b(n3270), .O(n3407));
  andx g3367(.a(n3203), .b(n345), .O(n3408));
  andx g3368(.a(n3408), .b(n3407), .O(n3409));
  andx g3369(.a(n3409), .b(n3405), .O(n3410));
  andx g3370(.a(n3359), .b(n922), .O(n3411));
  andx g3371(.a(n1942), .b(n3193), .O(n3412));
  andx g3372(.a(n3412), .b(n3298), .O(n3413));
  andx g3373(.a(n3413), .b(n3411), .O(n3414));
  orx  g3374(.a(n3414), .b(n3410), .O(n3415));
  andx g3375(.a(n107), .b(n75), .O(n3416));
  andx g3376(.a(n3416), .b(n42), .O(n3417));
  andx g3377(.a(n3417), .b(n431), .O(n3418));
  andx g3378(.a(n303), .b(n1687), .O(n3419));
  andx g3379(.a(n46), .b(n249), .O(n3420));
  andx g3380(.a(n3420), .b(n3419), .O(n3421));
  andx g3381(.a(n47), .b(pi35), .O(n3422));
  andx g3382(.a(n3422), .b(n1831), .O(n3423));
  andx g3383(.a(n3423), .b(n298), .O(n3424));
  andx g3384(.a(n3424), .b(n3421), .O(n3425));
  andx g3385(.a(n3425), .b(n3418), .O(n3426));
  andx g3386(.a(n3193), .b(n63), .O(n3427));
  andx g3387(.a(n42), .b(pi07), .O(n3428));
  andx g3388(.a(n3428), .b(n3240), .O(n3429));
  andx g3389(.a(n3429), .b(n3427), .O(n3430));
  andx g3390(.a(n3430), .b(n3394), .O(n3431));
  andx g3391(.a(n3246), .b(n67), .O(n3432));
  andx g3392(.a(n3203), .b(n430), .O(n3433));
  andx g3393(.a(n3433), .b(n3432), .O(n3434));
  andx g3394(.a(n3434), .b(n3431), .O(n3435));
  orx  g3395(.a(n3435), .b(n3426), .O(n3436));
  orx  g3396(.a(n3436), .b(n3415), .O(n3437));
  andx g3397(.a(n3383), .b(n313), .O(n3438));
  andx g3398(.a(n3438), .b(n3381), .O(n3439));
  andx g3399(.a(n3439), .b(n3361), .O(n3440));
  andx g3400(.a(n3344), .b(n93), .O(n3441));
  andx g3401(.a(n3340), .b(n3270), .O(n3442));
  andx g3402(.a(n3442), .b(n3441), .O(n3443));
  orx  g3403(.a(n3443), .b(n3440), .O(n3444));
  andx g3404(.a(n3253), .b(n67), .O(n3445));
  andx g3405(.a(n3445), .b(n3354), .O(n3446));
  andx g3406(.a(n3418), .b(n1831), .O(n3447));
  andx g3407(.a(n3447), .b(n3446), .O(n3448));
  andx g3408(.a(n3314), .b(n3195), .O(n3449));
  andx g3409(.a(n3449), .b(n644), .O(n3450));
  andx g3410(.a(n43), .b(pi35), .O(n3451));
  andx g3411(.a(n249), .b(n63), .O(n3452));
  andx g3412(.a(n3452), .b(n3451), .O(n3453));
  andx g3413(.a(n545), .b(n48), .O(n3454));
  andx g3414(.a(n3454), .b(n3453), .O(n3455));
  andx g3415(.a(n3455), .b(n3450), .O(n3456));
  orx  g3416(.a(n3456), .b(n3448), .O(n3457));
  orx  g3417(.a(n3457), .b(n3444), .O(n3458));
  orx  g3418(.a(n3458), .b(n3437), .O(n3459));
  orx  g3419(.a(n3459), .b(n3401), .O(n3460));
  orx  g3420(.a(n3460), .b(n3339), .O(n3461));
  andx g3421(.a(pi20), .b(n93), .O(n3462));
  andx g3422(.a(n3462), .b(pi17), .O(n3463));
  andx g3423(.a(n3463), .b(n3230), .O(n3464));
  andx g3424(.a(n3231), .b(n87), .O(n3465));
  andx g3425(.a(n3465), .b(n3386), .O(n3466));
  andx g3426(.a(n3466), .b(n3464), .O(n3467));
  andx g3427(.a(n48), .b(n63), .O(n3468));
  andx g3428(.a(pi35), .b(n67), .O(n3469));
  andx g3429(.a(n3469), .b(n3221), .O(n3470));
  andx g3430(.a(n3470), .b(n3468), .O(n3471));
  andx g3431(.a(n3471), .b(n3245), .O(n3472));
  orx  g3432(.a(n3472), .b(n3467), .O(n3473));
  andx g3433(.a(n3203), .b(n93), .O(n3474));
  andx g3434(.a(n3474), .b(n3359), .O(n3475));
  andx g3435(.a(n3290), .b(n87), .O(n3476));
  andx g3436(.a(n3218), .b(n3199), .O(n3477));
  andx g3437(.a(n3477), .b(n3476), .O(n3478));
  andx g3438(.a(n3478), .b(n3475), .O(n3479));
  andx g3439(.a(n3290), .b(n91), .O(n3480));
  andx g3440(.a(n3212), .b(n1021), .O(n3481));
  andx g3441(.a(n3481), .b(n3480), .O(n3482));
  andx g3442(.a(n3482), .b(n3269), .O(n3483));
  orx  g3443(.a(n3483), .b(n3479), .O(n3484));
  orx  g3444(.a(n3484), .b(n3473), .O(n3485));
  andx g3445(.a(n3394), .b(n3243), .O(n3486));
  andx g3446(.a(n3486), .b(n3250), .O(n3487));
  andx g3447(.a(n3267), .b(pi16), .O(n3488));
  andx g3448(.a(n3488), .b(pi20), .O(n3489));
  andx g3449(.a(n1942), .b(n91), .O(n3490));
  andx g3450(.a(n3490), .b(n3180), .O(n3491));
  andx g3451(.a(n3491), .b(n3489), .O(n3492));
  orx  g3452(.a(n3492), .b(n3487), .O(n3493));
  andx g3453(.a(n3406), .b(n1831), .O(n3494));
  andx g3454(.a(n3494), .b(n3203), .O(n3495));
  andx g3455(.a(n3214), .b(n1689), .O(n3496));
  andx g3456(.a(n3496), .b(n3495), .O(n3497));
  andx g3457(.a(n3497), .b(n3418), .O(n3498));
  andx g3458(.a(n3365), .b(n3259), .O(n3499));
  andx g3459(.a(n3406), .b(n164), .O(n3500));
  andx g3460(.a(n3382), .b(n3367), .O(n3501));
  andx g3461(.a(n3501), .b(n3500), .O(n3502));
  andx g3462(.a(n3502), .b(n3271), .O(n3503));
  andx g3463(.a(n3503), .b(n3499), .O(n3504));
  orx  g3464(.a(n3504), .b(n3498), .O(n3505));
  orx  g3465(.a(n3505), .b(n3493), .O(n3506));
  orx  g3466(.a(n3506), .b(n3485), .O(n3507));
  andx g3467(.a(n93), .b(pi35), .O(n3508));
  andx g3468(.a(n3508), .b(n45), .O(n3509));
  andx g3469(.a(n3509), .b(n3468), .O(n3510));
  andx g3470(.a(n3344), .b(n88), .O(n3511));
  andx g3471(.a(n3511), .b(n3510), .O(n3512));
  andx g3472(.a(n3305), .b(n449), .O(n3513));
  andx g3473(.a(n3513), .b(n3427), .O(n3514));
  andx g3474(.a(n3514), .b(n3796), .O(n3515));
  andx g3475(.a(n3508), .b(n3231), .O(n3516));
  andx g3476(.a(n3516), .b(n3515), .O(n3517));
  andx g3477(.a(pi16), .b(n3187), .O(n3518));
  andx g3478(.a(n3518), .b(pi20), .O(n3519));
  andx g3479(.a(n3285), .b(n3184), .O(n3520));
  andx g3480(.a(n3520), .b(n3519), .O(n3521));
  andx g3481(.a(n3521), .b(pi35), .O(n3522));
  andx g3482(.a(n3522), .b(n3328), .O(n3523));
  orx  g3483(.a(n3523), .b(n3517), .O(n3524));
  orx  g3484(.a(n3524), .b(n3512), .O(n3525));
  andx g3485(.a(n3402), .b(n329), .O(n3526));
  andx g3486(.a(n3526), .b(n64), .O(n3527));
  andx g3487(.a(n3527), .b(n3223), .O(n3528));
  andx g3488(.a(n93), .b(n212), .O(n3529));
  andx g3489(.a(n3529), .b(n64), .O(n3530));
  andx g3490(.a(n3530), .b(n3295), .O(n3531));
  andx g3491(.a(n3199), .b(n87), .O(n3532));
  andx g3492(.a(n3532), .b(n3354), .O(n3533));
  andx g3493(.a(n3533), .b(n3531), .O(n3534));
  orx  g3494(.a(n3534), .b(n3528), .O(n3535));
  andx g3495(.a(n3290), .b(n1503), .O(n3536));
  andx g3496(.a(n3536), .b(n2076), .O(n3537));
  andx g3497(.a(n3389), .b(pi18), .O(n3538));
  andx g3498(.a(n3538), .b(n3305), .O(n3539));
  andx g3499(.a(n93), .b(n3187), .O(n3540));
  andx g3500(.a(n3540), .b(n3539), .O(n3541));
  andx g3501(.a(n3541), .b(n3537), .O(n3542));
  andx g3502(.a(n3230), .b(n3189), .O(n3543));
  andx g3503(.a(n431), .b(n3193), .O(n3544));
  andx g3504(.a(n3469), .b(n92), .O(n3545));
  andx g3505(.a(n3545), .b(n3544), .O(n3546));
  andx g3506(.a(n3546), .b(n3543), .O(n3547));
  orx  g3507(.a(n3547), .b(n3542), .O(n3548));
  orx  g3508(.a(n3548), .b(n3535), .O(n3549));
  orx  g3509(.a(n3549), .b(n3525), .O(n3550));
  orx  g3510(.a(n3550), .b(n3507), .O(n3551));
  andx g3511(.a(n3427), .b(n107), .O(n3552));
  andx g3512(.a(n2682), .b(n64), .O(n3553));
  andx g3513(.a(n3553), .b(n2256), .O(n3554));
  andx g3514(.a(n3554), .b(n3552), .O(n3555));
  andx g3515(.a(n46), .b(pi09), .O(n3556));
  andx g3516(.a(n3556), .b(n67), .O(n3557));
  andx g3517(.a(n3557), .b(n3354), .O(n3558));
  andx g3518(.a(n3558), .b(n3555), .O(n3559));
  andx g3519(.a(n3268), .b(n3190), .O(n3560));
  andx g3520(.a(n3560), .b(n3491), .O(n3561));
  orx  g3521(.a(n3561), .b(n3559), .O(n3562));
  andx g3522(.a(n3320), .b(n3193), .O(n3563));
  andx g3523(.a(pi35), .b(n87), .O(n3564));
  andx g3524(.a(n3564), .b(n895), .O(n3565));
  andx g3525(.a(n3565), .b(n3563), .O(n3566));
  andx g3526(.a(n3306), .b(n3184), .O(n3567));
  andx g3527(.a(n3567), .b(n3188), .O(n3568));
  andx g3528(.a(n3568), .b(n3566), .O(n3569));
  andx g3529(.a(n3346), .b(n48), .O(n3570));
  andx g3530(.a(n3570), .b(n3453), .O(n3571));
  andx g3531(.a(n3571), .b(n3441), .O(n3572));
  orx  g3532(.a(n3572), .b(n3569), .O(n3573));
  orx  g3533(.a(n3573), .b(n3562), .O(n3574));
  andx g3534(.a(n3270), .b(n67), .O(n3575));
  andx g3535(.a(n3575), .b(n3222), .O(n3576));
  andx g3536(.a(n42), .b(n75), .O(n3577));
  andx g3537(.a(n3577), .b(n3552), .O(n3578));
  andx g3538(.a(n73), .b(n533), .O(n3579));
  andx g3539(.a(n3579), .b(n3578), .O(n3580));
  andx g3540(.a(n3580), .b(n3576), .O(n3581));
  andx g3541(.a(n3242), .b(n431), .O(n3582));
  andx g3542(.a(n3582), .b(n3244), .O(n3583));
  andx g3543(.a(n3583), .b(n3304), .O(n3584));
  orx  g3544(.a(n3584), .b(n3581), .O(n3585));
  andx g3545(.a(n3298), .b(n3563), .O(n3586));
  andx g3546(.a(n3586), .b(n3464), .O(n3587));
  andx g3547(.a(n1758), .b(n48), .O(n3588));
  andx g3548(.a(n3202), .b(n164), .O(n3589));
  andx g3549(.a(n3589), .b(n45), .O(n3590));
  andx g3550(.a(n3590), .b(n3588), .O(n3591));
  andx g3551(.a(n3591), .b(n3366), .O(n3592));
  orx  g3552(.a(n3592), .b(n3587), .O(n3593));
  orx  g3553(.a(n3593), .b(n3585), .O(n3594));
  orx  g3554(.a(n3594), .b(n3574), .O(n3595));
  andx g3555(.a(n3533), .b(n3450), .O(n3596));
  andx g3556(.a(n3297), .b(n3214), .O(n3597));
  andx g3557(.a(n3597), .b(n3272), .O(n3598));
  andx g3558(.a(n3598), .b(n3321), .O(n3599));
  andx g3559(.a(n3599), .b(n3319), .O(n3600));
  orx  g3560(.a(n3600), .b(n3596), .O(n3601));
  andx g3561(.a(n2832), .b(n48), .O(n3602));
  andx g3562(.a(n3602), .b(n3280), .O(n3603));
  andx g3563(.a(n3603), .b(n3279), .O(n3604));
  andx g3564(.a(n48), .b(pi35), .O(n3605));
  andx g3565(.a(n164), .b(n45), .O(n3606));
  andx g3566(.a(n3606), .b(n3605), .O(n3607));
  andx g3567(.a(n3194), .b(n431), .O(n3608));
  andx g3568(.a(n3608), .b(n42), .O(n3609));
  andx g3569(.a(n3609), .b(n41), .O(n3610));
  andx g3570(.a(n3610), .b(n3607), .O(n3611));
  orx  g3571(.a(n3611), .b(n3604), .O(n3612));
  orx  g3572(.a(n3612), .b(n3601), .O(n3613));
  andx g3573(.a(n3449), .b(n73), .O(n3614));
  andx g3574(.a(n3614), .b(n3510), .O(n3615));
  andx g3575(.a(n3232), .b(n855), .O(n3616));
  andx g3576(.a(n3616), .b(n3181), .O(n3617));
  andx g3577(.a(n3617), .b(n3522), .O(n3618));
  orx  g3578(.a(n3618), .b(n3615), .O(n3619));
  andx g3579(.a(n3214), .b(n1768), .O(n3620));
  andx g3580(.a(n3620), .b(n3393), .O(n3621));
  andx g3581(.a(n3621), .b(n3568), .O(n3622));
  andx g3582(.a(n3406), .b(n357), .O(n3623));
  andx g3583(.a(n41), .b(pi35), .O(n3624));
  andx g3584(.a(n3624), .b(n3203), .O(n3625));
  andx g3585(.a(n3625), .b(n3623), .O(n3626));
  andx g3586(.a(n3626), .b(n3405), .O(n3627));
  orx  g3587(.a(n3627), .b(n3622), .O(n3628));
  orx  g3588(.a(n3628), .b(n3619), .O(n3629));
  orx  g3589(.a(n3629), .b(n3613), .O(n3630));
  orx  g3590(.a(n3630), .b(n3595), .O(n3631));
  orx  g3591(.a(n3631), .b(n3551), .O(n3632));
  orx  g3592(.a(n3632), .b(n3461), .O(n3633));
  andx g3593(.a(n3529), .b(n3203), .O(n3634));
  andx g3594(.a(n3634), .b(n3381), .O(n3635));
  andx g3595(.a(n3297), .b(n3193), .O(n3636));
  andx g3596(.a(n3270), .b(n3199), .O(n3637));
  andx g3597(.a(n3637), .b(n3636), .O(n3638));
  andx g3598(.a(n3638), .b(n3635), .O(n3639));
  andx g3599(.a(n3469), .b(n3340), .O(n3640));
  andx g3600(.a(n3194), .b(n60), .O(n3641));
  andx g3601(.a(pi16), .b(pi15), .O(n3642));
  andx g3602(.a(n3642), .b(n3641), .O(n3643));
  andx g3603(.a(pi07), .b(pi19), .O(n3644));
  andx g3604(.a(n3644), .b(n64), .O(n3645));
  andx g3605(.a(n3645), .b(n3643), .O(n3646));
  andx g3606(.a(n3646), .b(n3640), .O(n3647));
  orx  g3607(.a(n3647), .b(n3639), .O(n3648));
  andx g3608(.a(n303), .b(n212), .O(n3649));
  andx g3609(.a(n3649), .b(n3367), .O(n3650));
  andx g3610(.a(n3650), .b(n3370), .O(n3651));
  andx g3611(.a(n3651), .b(n3271), .O(n3652));
  andx g3612(.a(n3652), .b(n3499), .O(n3653));
  andx g3613(.a(n3295), .b(n3262), .O(n3654));
  andx g3614(.a(n3654), .b(n3356), .O(n3655));
  orx  g3615(.a(n3655), .b(n3653), .O(n3656));
  orx  g3616(.a(n3656), .b(n3648), .O(n3657));
  andx g3617(.a(n3427), .b(n250), .O(n3658));
  andx g3618(.a(n3565), .b(n3189), .O(n3659));
  andx g3619(.a(n3659), .b(n3658), .O(n3660));
  andx g3620(.a(n3660), .b(n3230), .O(n3661));
  andx g3621(.a(n3185), .b(pi16), .O(n3662));
  andx g3622(.a(n3662), .b(pi20), .O(n3663));
  andx g3623(.a(n3215), .b(n313), .O(n3664));
  andx g3624(.a(n3664), .b(n3663), .O(n3665));
  orx  g3625(.a(n3665), .b(n3661), .O(n3666));
  andx g3626(.a(n48), .b(pi09), .O(n3667));
  andx g3627(.a(n3667), .b(n3509), .O(n3668));
  andx g3628(.a(n3668), .b(n3555), .O(n3669));
  andx g3629(.a(n3389), .b(n3365), .O(n3670));
  andx g3630(.a(n3253), .b(n63), .O(n3671));
  andx g3631(.a(n533), .b(pi35), .O(n3672));
  andx g3632(.a(n3672), .b(n3203), .O(n3673));
  andx g3633(.a(n3673), .b(n313), .O(n3674));
  andx g3634(.a(n3674), .b(n3671), .O(n3675));
  andx g3635(.a(n3675), .b(n3670), .O(n3676));
  orx  g3636(.a(n3676), .b(n3669), .O(n3677));
  orx  g3637(.a(n3677), .b(n3666), .O(n3678));
  orx  g3638(.a(n3678), .b(n3657), .O(n3679));
  andx g3639(.a(n3417), .b(n3239), .O(n3680));
  andx g3640(.a(n3234), .b(n1689), .O(n3681));
  andx g3641(.a(n3681), .b(n3495), .O(n3682));
  andx g3642(.a(n3682), .b(n3680), .O(n3683));
  andx g3643(.a(n1344), .b(n60), .O(n3684));
  andx g3644(.a(n3684), .b(n333), .O(n3685));
  andx g3645(.a(n3685), .b(n3519), .O(n3686));
  andx g3646(.a(n3214), .b(n63), .O(n3687));
  andx g3647(.a(n3687), .b(n3273), .O(n3688));
  andx g3648(.a(n3688), .b(n3686), .O(n3689));
  orx  g3649(.a(n3689), .b(n3683), .O(n3690));
  andx g3650(.a(n3451), .b(n3261), .O(n3691));
  andx g3651(.a(n3691), .b(n313), .O(n3692));
  andx g3652(.a(n3692), .b(n3588), .O(n3693));
  andx g3653(.a(n3693), .b(n3499), .O(n3694));
  andx g3654(.a(n3518), .b(n3285), .O(n3695));
  andx g3655(.a(n3695), .b(n3194), .O(n3696));
  andx g3656(.a(n3696), .b(n73), .O(n3697));
  andx g3657(.a(n3234), .b(n91), .O(n3698));
  andx g3658(.a(n3698), .b(n3248), .O(n3699));
  andx g3659(.a(n3699), .b(n3697), .O(n3700));
  orx  g3660(.a(n3700), .b(n3694), .O(n3701));
  orx  g3661(.a(n3701), .b(n3690), .O(n3702));
  andx g3662(.a(n3582), .b(n3394), .O(n3703));
  andx g3663(.a(n3703), .b(n3304), .O(n3704));
  andx g3664(.a(n1344), .b(pi16), .O(n3705));
  andx g3665(.a(n3705), .b(n3389), .O(n3706));
  andx g3666(.a(n3706), .b(n43), .O(n3707));
  andx g3667(.a(n533), .b(n47), .O(n3708));
  andx g3668(.a(n2832), .b(n895), .O(n3709));
  andx g3669(.a(n3709), .b(n3708), .O(n3710));
  andx g3670(.a(n3710), .b(n3247), .O(n3711));
  andx g3671(.a(n3711), .b(n3707), .O(n3712));
  orx  g3672(.a(n3712), .b(n3704), .O(n3713));
  andx g3673(.a(n3258), .b(n3196), .O(n3714));
  andx g3674(.a(n3714), .b(n3352), .O(n3715));
  andx g3675(.a(n3715), .b(n3446), .O(n3716));
  andx g3676(.a(n3365), .b(n3314), .O(n3717));
  andx g3677(.a(n3234), .b(n895), .O(n3718));
  andx g3678(.a(n43), .b(n64), .O(n3719));
  andx g3679(.a(n3719), .b(n3218), .O(n3720));
  andx g3680(.a(n3720), .b(n48), .O(n3721));
  andx g3681(.a(n3721), .b(n3718), .O(n3722));
  andx g3682(.a(n3722), .b(n3717), .O(n3723));
  orx  g3683(.a(n3723), .b(n3716), .O(n3724));
  orx  g3684(.a(n3724), .b(n3713), .O(n3725));
  orx  g3685(.a(n3725), .b(n3702), .O(n3726));
  orx  g3686(.a(n3726), .b(n3679), .O(n3727));
  andx g3687(.a(n3469), .b(n49), .O(n3728));
  andx g3688(.a(n3728), .b(n1810), .O(n3729));
  andx g3689(.a(n3729), .b(n3449), .O(n3730));
  andx g3690(.a(n60), .b(n42), .O(n3731));
  andx g3691(.a(n3731), .b(n3390), .O(n3732));
  andx g3692(.a(n3732), .b(n88), .O(n3733));
  andx g3693(.a(n3422), .b(n3369), .O(n3734));
  andx g3694(.a(pi19), .b(n64), .O(n3735));
  andx g3695(.a(n3187), .b(n63), .O(n3736));
  andx g3696(.a(n3736), .b(n3735), .O(n3737));
  andx g3697(.a(n3737), .b(n3734), .O(n3738));
  andx g3698(.a(n3738), .b(n3385), .O(n3739));
  andx g3699(.a(n3739), .b(n3733), .O(n3740));
  orx  g3700(.a(n3740), .b(n3730), .O(n3741));
  andx g3701(.a(n3706), .b(n93), .O(n3742));
  andx g3702(.a(n3708), .b(n3219), .O(n3743));
  andx g3703(.a(n3743), .b(n3221), .O(n3744));
  andx g3704(.a(n3744), .b(n3671), .O(n3745));
  andx g3705(.a(n3745), .b(n3742), .O(n3746));
  andx g3706(.a(n3197), .b(n43), .O(n3747));
  andx g3707(.a(n855), .b(n557), .O(n3748));
  andx g3708(.a(n3202), .b(n644), .O(n3749));
  andx g3709(.a(n3749), .b(n48), .O(n3750));
  andx g3710(.a(n3750), .b(n3748), .O(n3751));
  andx g3711(.a(n3751), .b(n3747), .O(n3752));
  orx  g3712(.a(n3752), .b(n3746), .O(n3753));
  orx  g3713(.a(n3753), .b(n3741), .O(n3754));
  andx g3714(.a(n3290), .b(n93), .O(n3755));
  andx g3715(.a(n3212), .b(n3181), .O(n3756));
  andx g3716(.a(n3756), .b(n3755), .O(n3757));
  andx g3717(.a(n3757), .b(n3686), .O(n3758));
  andx g3718(.a(n3218), .b(n303), .O(n3759));
  andx g3719(.a(n46), .b(pi07), .O(n3760));
  andx g3720(.a(n3760), .b(n3255), .O(n3761));
  andx g3721(.a(n3761), .b(n3691), .O(n3762));
  andx g3722(.a(n3762), .b(n3759), .O(n3763));
  andx g3723(.a(n3763), .b(n3260), .O(n3764));
  orx  g3724(.a(n3764), .b(n3758), .O(n3765));
  andx g3725(.a(n3367), .b(n545), .O(n3766));
  andx g3726(.a(n3369), .b(n3261), .O(n3767));
  andx g3727(.a(n3767), .b(n3766), .O(n3768));
  andx g3728(.a(n3768), .b(n3575), .O(n3769));
  andx g3729(.a(n3769), .b(n3260), .O(n3770));
  andx g3730(.a(n3318), .b(n3286), .O(n3771));
  andx g3731(.a(pi20), .b(n67), .O(n3772));
  andx g3732(.a(n3772), .b(n3597), .O(n3773));
  andx g3733(.a(n3773), .b(n3321), .O(n3774));
  andx g3734(.a(n3774), .b(n3771), .O(n3775));
  orx  g3735(.a(n3775), .b(n3770), .O(n3776));
  orx  g3736(.a(n3776), .b(n3765), .O(n3777));
  orx  g3737(.a(n3777), .b(n3754), .O(n3778));
  andx g3738(.a(n3511), .b(n3356), .O(n3779));
  andx g3739(.a(n3719), .b(n313), .O(n3780));
  andx g3740(.a(n3780), .b(n3605), .O(n3781));
  andx g3741(.a(n3781), .b(n3610), .O(n3782));
  orx  g3742(.a(n3782), .b(n3779), .O(n3783));
  andx g3743(.a(n3234), .b(n3193), .O(n3784));
  andx g3744(.a(n3413), .b(n3384), .O(n3785));
  andx g3745(.a(pi18), .b(pi16), .O(n3786));
  andx g3746(.a(n3786), .b(n42), .O(n3787));
  andx g3747(.a(n3787), .b(n3208), .O(n3788));
  andx g3748(.a(n431), .b(n333), .O(n3789));
  andx g3749(.a(n3248), .b(n1454), .O(n3790));
  andx g3750(.a(n3790), .b(n3214), .O(n3791));
  andx g3751(.a(n3791), .b(n3789), .O(n3792));
  andx g3752(.a(n3792), .b(n3788), .O(n3793));
  orx  g3753(.a(n3793), .b(n3785), .O(n3794));
  orx  g3754(.a(n3794), .b(n3783), .O(n3795));
  andx g3755(.a(n3644), .b(n3187), .O(n3796));
  andx g3756(.a(n3796), .b(n345), .O(n3797));
  andx g3757(.a(n3797), .b(n3307), .O(n3798));
  andx g3758(.a(n3798), .b(n3304), .O(n3799));
  andx g3759(.a(n3614), .b(n3356), .O(n3800));
  orx  g3760(.a(n3800), .b(n3799), .O(n3801));
  andx g3761(.a(n3180), .b(n63), .O(n3802));
  andx g3762(.a(n3272), .b(n3181), .O(n3803));
  andx g3763(.a(n3803), .b(n3802), .O(n3804));
  andx g3764(.a(n3804), .b(n3211), .O(n3805));
  andx g3765(.a(n3290), .b(n1901), .O(n3806));
  andx g3766(.a(n3806), .b(n3515), .O(n3807));
  orx  g3767(.a(n3807), .b(n3805), .O(n3808));
  orx  g3768(.a(n3808), .b(n3801), .O(n3809));
  orx  g3769(.a(n3809), .b(n3795), .O(n3810));
  orx  g3770(.a(n3810), .b(n3778), .O(n3811));
  orx  g3771(.a(n3811), .b(n3727), .O(n3812));
  andx g3772(.a(n3341), .b(n45), .O(n3813));
  andx g3773(.a(n3813), .b(n3468), .O(n3814));
  andx g3774(.a(n3814), .b(n3717), .O(n3815));
  andx g3775(.a(n3513), .b(n3320), .O(n3816));
  andx g3776(.a(n3816), .b(n3796), .O(n3817));
  andx g3777(.a(n3248), .b(n3214), .O(n3818));
  andx g3778(.a(n3818), .b(n3817), .O(n3819));
  orx  g3779(.a(n3819), .b(n3815), .O(n3820));
  andx g3780(.a(pi35), .b(n3193), .O(n3821));
  andx g3781(.a(n3821), .b(n431), .O(n3822));
  andx g3782(.a(n3822), .b(n3360), .O(n3823));
  andx g3783(.a(n3680), .b(n1831), .O(n3824));
  andx g3784(.a(n3824), .b(n3510), .O(n3825));
  orx  g3785(.a(n3825), .b(n3823), .O(n3826));
  orx  g3786(.a(n3826), .b(n3820), .O(n3827));
  andx g3787(.a(n3297), .b(n3234), .O(n3828));
  andx g3788(.a(n3719), .b(n3348), .O(n3829));
  andx g3789(.a(n3829), .b(n3828), .O(n3830));
  andx g3790(.a(n3830), .b(n3449), .O(n3831));
  andx g3791(.a(n3231), .b(n75), .O(n3832));
  andx g3792(.a(n3736), .b(n3232), .O(n3833));
  andx g3793(.a(n3833), .b(n3214), .O(n3834));
  andx g3794(.a(n3834), .b(n3832), .O(n3835));
  andx g3795(.a(n3835), .b(n3539), .O(n3836));
  orx  g3796(.a(n3836), .b(n3831), .O(n3837));
  andx g3797(.a(n3221), .b(n73), .O(n3838));
  andx g3798(.a(n3838), .b(n3214), .O(n3839));
  andx g3799(.a(n3839), .b(n3348), .O(n3840));
  andx g3800(.a(n3840), .b(n3315), .O(n3841));
  andx g3801(.a(n3643), .b(n64), .O(n3842));
  andx g3802(.a(n1901), .b(n87), .O(n3843));
  andx g3803(.a(n3290), .b(n3212), .O(n3844));
  andx g3804(.a(n3844), .b(n3843), .O(n3845));
  andx g3805(.a(n3845), .b(n3842), .O(n3846));
  orx  g3806(.a(n3846), .b(n3841), .O(n3847));
  orx  g3807(.a(n3847), .b(n3837), .O(n3848));
  orx  g3808(.a(n3848), .b(n3827), .O(n3849));
  andx g3809(.a(n3209), .b(n3194), .O(n3850));
  andx g3810(.a(n3850), .b(n3189), .O(n3851));
  andx g3811(.a(n1503), .b(pi35), .O(n3852));
  andx g3812(.a(n3852), .b(n3213), .O(n3853));
  andx g3813(.a(n3853), .b(n3851), .O(n3854));
  andx g3814(.a(pi35), .b(n91), .O(n3855));
  andx g3815(.a(n533), .b(n63), .O(n3856));
  andx g3816(.a(n3856), .b(n3297), .O(n3857));
  andx g3817(.a(n3857), .b(n3855), .O(n3858));
  andx g3818(.a(n3858), .b(n3392), .O(n3859));
  orx  g3819(.a(n3859), .b(n3854), .O(n3860));
  andx g3820(.a(n3287), .b(n64), .O(n3861));
  andx g3821(.a(n3861), .b(n3566), .O(n3862));
  andx g3822(.a(n3446), .b(n3316), .O(n3863));
  orx  g3823(.a(n3863), .b(n3862), .O(n3864));
  orx  g3824(.a(n3864), .b(n3860), .O(n3865));
  andx g3825(.a(n3344), .b(n41), .O(n3866));
  andx g3826(.a(n3866), .b(n3510), .O(n3867));
  andx g3827(.a(n3866), .b(n3356), .O(n3868));
  orx  g3828(.a(n3868), .b(n3867), .O(n3869));
  andx g3829(.a(n3419), .b(n3270), .O(n3870));
  andx g3830(.a(n46), .b(n41), .O(n3871));
  andx g3831(.a(n2508), .b(n3870), .O(n3872));
  andx g3832(.a(n3872), .b(n3225), .O(n3873));
  andx g3833(.a(n3861), .b(n3621), .O(n3874));
  orx  g3834(.a(n3874), .b(n3873), .O(n3875));
  orx  g3835(.a(n3875), .b(n3869), .O(n3876));
  orx  g3836(.a(n3876), .b(n3865), .O(n3877));
  orx  g3837(.a(n3877), .b(n3849), .O(n3878));
  andx g3838(.a(n3429), .b(n855), .O(n3879));
  andx g3839(.a(n3246), .b(n93), .O(n3880));
  andx g3840(.a(n43), .b(n1687), .O(n3881));
  andx g3841(.a(n3881), .b(n3708), .O(n3882));
  andx g3842(.a(n3882), .b(n345), .O(n3883));
  andx g3843(.a(n3883), .b(n3880), .O(n3884));
  andx g3844(.a(n3884), .b(n3879), .O(n3885));
  andx g3845(.a(n3391), .b(n43), .O(n3886));
  andx g3846(.a(n3708), .b(n3199), .O(n3887));
  andx g3847(.a(n3887), .b(n3219), .O(n3888));
  andx g3848(.a(n3888), .b(n3385), .O(n3889));
  andx g3849(.a(n3889), .b(n3886), .O(n3890));
  orx  g3850(.a(n3890), .b(n3885), .O(n3891));
  andx g3851(.a(n3822), .b(n3439), .O(n3892));
  andx g3852(.a(n3771), .b(n3462), .O(n3893));
  andx g3853(.a(n3893), .b(n3537), .O(n3894));
  orx  g3854(.a(n3894), .b(n3892), .O(n3895));
  orx  g3855(.a(n3895), .b(n3891), .O(n3896));
  andx g3856(.a(n3358), .b(n3196), .O(n3897));
  andx g3857(.a(n46), .b(pi14), .O(n3898));
  andx g3858(.a(n3898), .b(n47), .O(n3899));
  andx g3859(.a(n3899), .b(n45), .O(n3900));
  andx g3860(.a(n3900), .b(n3897), .O(n3901));
  andx g3861(.a(n3784), .b(n3232), .O(n3902));
  andx g3862(.a(n3902), .b(n3901), .O(n3903));
  andx g3863(.a(n756), .b(pi14), .O(n3904));
  andx g3864(.a(n3904), .b(n3196), .O(n3905));
  andx g3865(.a(n3905), .b(n3552), .O(n3906));
  andx g3866(.a(n3906), .b(n3668), .O(n3907));
  orx  g3867(.a(n3907), .b(n3903), .O(n3908));
  andx g3868(.a(n3411), .b(n3387), .O(n3909));
  andx g3869(.a(n44), .b(n46), .O(n3910));
  andx g3870(.a(n93), .b(pi14), .O(n3911));
  andx g3871(.a(n3911), .b(n49), .O(n3912));
  andx g3872(.a(n3912), .b(n3897), .O(n3913));
  andx g3873(.a(n3913), .b(n3361), .O(n3914));
  orx  g3874(.a(n3914), .b(n3909), .O(n3915));
  orx  g3875(.a(n3915), .b(n3908), .O(n3916));
  orx  g3876(.a(n3916), .b(n3896), .O(n3917));
  andx g3877(.a(n3772), .b(n3239), .O(n3918));
  andx g3878(.a(n3918), .b(n3290), .O(n3919));
  andx g3879(.a(n3919), .b(n3321), .O(n3920));
  andx g3880(.a(n3920), .b(n3771), .O(n3921));
  andx g3881(.a(n895), .b(n249), .O(n3922));
  andx g3882(.a(n3369), .b(n73), .O(n3923));
  andx g3883(.a(n3923), .b(n3368), .O(n3924));
  andx g3884(.a(n3924), .b(n3922), .O(n3925));
  andx g3885(.a(n3925), .b(n3714), .O(n3926));
  orx  g3886(.a(n3926), .b(n3921), .O(n3927));
  andx g3887(.a(n3617), .b(n3332), .O(n3928));
  andx g3888(.a(n3455), .b(n3531), .O(n3929));
  orx  g3889(.a(n3929), .b(n3928), .O(n3930));
  orx  g3890(.a(n3930), .b(n3927), .O(n3931));
  andx g3891(.a(n3641), .b(n333), .O(n3932));
  andx g3892(.a(n3932), .b(n3519), .O(n3933));
  andx g3893(.a(n3508), .b(n3212), .O(n3934));
  andx g3894(.a(n3934), .b(n3465), .O(n3935));
  andx g3895(.a(n3935), .b(n3933), .O(n3936));
  andx g3896(.a(n533), .b(pi07), .O(n3937));
  andx g3897(.a(n3937), .b(n3578), .O(n3938));
  andx g3898(.a(n3938), .b(n3607), .O(n3939));
  orx  g3899(.a(n3939), .b(n3936), .O(n3940));
  andx g3900(.a(n3719), .b(n3202), .O(n3941));
  andx g3901(.a(n3941), .b(n313), .O(n3942));
  andx g3902(.a(n3942), .b(n3588), .O(n3943));
  andx g3903(.a(n3943), .b(n3366), .O(n3944));
  andx g3904(.a(n3699), .b(n3646), .O(n3945));
  orx  g3905(.a(n3945), .b(n3944), .O(n3946));
  orx  g3906(.a(n3946), .b(n3940), .O(n3947));
  orx  g3907(.a(n3947), .b(n3931), .O(n3948));
  orx  g3908(.a(n3948), .b(n3917), .O(n3949));
  orx  g3909(.a(n3949), .b(n3878), .O(n3950));
  orx  g3910(.a(n3950), .b(n3812), .O(n3951));
  orx  g3911(.a(n3951), .b(n3633), .O(n3952));
  andx g3912(.a(n46), .b(n3193), .O(n3953));
  andx g3913(.a(n3953), .b(n3290), .O(n3954));
  andx g3914(.a(n3954), .b(n230), .O(n3955));
  andx g3915(.a(n3788), .b(n41), .O(n3956));
  andx g3916(.a(n3956), .b(n3203), .O(n3957));
  andx g3917(.a(n3957), .b(n644), .O(n3958));
  andx g3918(.a(n3958), .b(n3955), .O(n3959));
  andx g3919(.a(n3788), .b(n88), .O(n3960));
  andx g3920(.a(n3960), .b(n3203), .O(n3961));
  andx g3921(.a(n3961), .b(n644), .O(n3962));
  andx g3922(.a(n3962), .b(n3955), .O(n3963));
  orx  g3923(.a(n3963), .b(n3959), .O(n3964));
  andx g3924(.a(n3234), .b(n67), .O(n3965));
  andx g3925(.a(n3965), .b(n3419), .O(n3966));
  andx g3926(.a(n3577), .b(pi18), .O(n3967));
  andx g3927(.a(n3967), .b(n3305), .O(n3968));
  andx g3928(.a(n3968), .b(n88), .O(n3969));
  andx g3929(.a(n3969), .b(n43), .O(n3970));
  andx g3930(.a(n46), .b(n3187), .O(n3971));
  andx g3931(.a(n3971), .b(n47), .O(n3972));
  andx g3932(.a(n3972), .b(n73), .O(n3973));
  andx g3933(.a(n3973), .b(n3970), .O(n3974));
  andx g3934(.a(n3974), .b(n3966), .O(n3975));
  andx g3935(.a(n855), .b(n3193), .O(n3976));
  andx g3936(.a(n3976), .b(n3469), .O(n3977));
  andx g3937(.a(n3977), .b(n3974), .O(n3978));
  orx  g3938(.a(n3978), .b(n3975), .O(n3979));
  orx  g3939(.a(n3979), .b(n3964), .O(n3980));
  andx g3940(.a(n3968), .b(n3187), .O(n3981));
  andx g3941(.a(n3981), .b(n43), .O(n3982));
  andx g3942(.a(n3871), .b(n47), .O(n3983));
  andx g3943(.a(n3983), .b(n644), .O(n3984));
  andx g3944(.a(n3984), .b(n3982), .O(n3985));
  andx g3945(.a(n3564), .b(n63), .O(n3986));
  andx g3946(.a(n3986), .b(n3419), .O(n3987));
  andx g3947(.a(n3987), .b(n3985), .O(n3988));
  andx g3948(.a(n3565), .b(n2076), .O(n3989));
  andx g3949(.a(n3960), .b(n922), .O(n3990));
  andx g3950(.a(n3990), .b(n64), .O(n3991));
  andx g3951(.a(n3991), .b(n3989), .O(n3992));
  orx  g3952(.a(n3992), .b(n3988), .O(n3993));
  andx g3953(.a(n3306), .b(n3284), .O(n3994));
  andx g3954(.a(n3994), .b(n41), .O(n3995));
  andx g3955(.a(n3995), .b(n43), .O(n3996));
  andx g3956(.a(n3760), .b(n47), .O(n3997));
  andx g3957(.a(n3997), .b(n3735), .O(n3998));
  andx g3958(.a(n3998), .b(n3996), .O(n3999));
  andx g3959(.a(n3999), .b(n3977), .O(n4000));
  andx g3960(.a(n1344), .b(n333), .O(n4001));
  andx g3961(.a(n3821), .b(n855), .O(n4002));
  andx g3962(.a(n4002), .b(n4001), .O(n4003));
  andx g3963(.a(n3990), .b(n93), .O(n4004));
  andx g3964(.a(n4004), .b(n4003), .O(n4005));
  orx  g3965(.a(n4005), .b(n4000), .O(n4006));
  orx  g3966(.a(n4006), .b(n3993), .O(n4007));
  orx  g3967(.a(n4007), .b(n3980), .O(n4008));
  andx g3968(.a(n3961), .b(n73), .O(n4009));
  andx g3969(.a(n3214), .b(n3199), .O(n4010));
  andx g3970(.a(n895), .b(n75), .O(n4011));
  andx g3971(.a(n4011), .b(n4010), .O(n4012));
  andx g3972(.a(n4012), .b(n4009), .O(n4013));
  andx g3973(.a(n3636), .b(n3234), .O(n4014));
  andx g3974(.a(n4014), .b(n3985), .O(n4015));
  orx  g3975(.a(n4015), .b(n4013), .O(n4016));
  andx g3976(.a(n3290), .b(n1758), .O(n4017));
  andx g3977(.a(n4017), .b(n4001), .O(n4018));
  andx g3978(.a(n4018), .b(n4004), .O(n4019));
  andx g3979(.a(n3983), .b(n73), .O(n4020));
  andx g3980(.a(n4020), .b(n3982), .O(n4021));
  andx g3981(.a(n4021), .b(n3966), .O(n4022));
  orx  g3982(.a(n4022), .b(n4019), .O(n4023));
  orx  g3983(.a(n4023), .b(n4016), .O(n4024));
  andx g3984(.a(n3994), .b(n88), .O(n4025));
  andx g3985(.a(n4025), .b(n43), .O(n4026));
  andx g3986(.a(n4026), .b(n3998), .O(n4027));
  andx g3987(.a(n4027), .b(n3977), .O(n4028));
  andx g3988(.a(n3297), .b(n75), .O(n4029));
  andx g3989(.a(n4029), .b(n4010), .O(n4030));
  andx g3990(.a(n4030), .b(n3958), .O(n4031));
  orx  g3991(.a(n4031), .b(n4028), .O(n4032));
  andx g3992(.a(n46), .b(pi19), .O(n4033));
  andx g3993(.a(n4033), .b(n47), .O(n4034));
  andx g3994(.a(n4034), .b(n644), .O(n4035));
  andx g3995(.a(n4035), .b(n3996), .O(n4036));
  andx g3996(.a(n4036), .b(n3987), .O(n4037));
  andx g3997(.a(n3821), .b(n895), .O(n4038));
  andx g3998(.a(n4038), .b(n230), .O(n4039));
  andx g3999(.a(n4039), .b(n3991), .O(n4040));
  orx  g4000(.a(n4040), .b(n4037), .O(n4041));
  orx  g4001(.a(n4041), .b(n4032), .O(n4042));
  orx  g4002(.a(n4042), .b(n4024), .O(n4043));
  orx  g4003(.a(n4043), .b(n4008), .O(n4044));
  andx g4004(.a(n3957), .b(n73), .O(n4045));
  andx g4005(.a(n3954), .b(n3402), .O(n4046));
  andx g4006(.a(n4046), .b(n4045), .O(n4047));
  andx g4007(.a(n3956), .b(n922), .O(n4048));
  andx g4008(.a(n4048), .b(n64), .O(n4049));
  andx g4009(.a(n3989), .b(n4049), .O(n4050));
  orx  g4010(.a(n4050), .b(n4047), .O(n4051));
  andx g4011(.a(n4046), .b(n4009), .O(n4052));
  andx g4012(.a(n4030), .b(n3962), .O(n4053));
  orx  g4013(.a(n4053), .b(n4052), .O(n4054));
  orx  g4014(.a(n4054), .b(n4051), .O(n4055));
  andx g4015(.a(n4048), .b(n93), .O(n4056));
  andx g4016(.a(n229), .b(n333), .O(n4057));
  andx g4017(.a(n4018), .b(n4056), .O(n4058));
  andx g4018(.a(n4049), .b(n4039), .O(n4059));
  orx  g4019(.a(n4059), .b(n4058), .O(n4060));
  andx g4020(.a(n4036), .b(n4014), .O(n4061));
  andx g4021(.a(n3972), .b(n644), .O(n4062));
  andx g4022(.a(n4062), .b(n3970), .O(n4063));
  andx g4023(.a(n4063), .b(n4014), .O(n4064));
  orx  g4024(.a(n4064), .b(n4061), .O(n4065));
  orx  g4025(.a(n4065), .b(n4060), .O(n4066));
  orx  g4026(.a(n4066), .b(n4055), .O(n4067));
  andx g4027(.a(n4035), .b(n4026), .O(n4068));
  andx g4028(.a(n4068), .b(n3987), .O(n4069));
  andx g4029(.a(n4027), .b(n3966), .O(n4070));
  orx  g4030(.a(n4070), .b(n4069), .O(n4071));
  andx g4031(.a(n3999), .b(n3966), .O(n4072));
  andx g4032(.a(n4068), .b(n4014), .O(n4073));
  orx  g4033(.a(n4073), .b(n4072), .O(n4074));
  orx  g4034(.a(n4074), .b(n4071), .O(n4075));
  andx g4035(.a(n4045), .b(n4012), .O(n4076));
  andx g4036(.a(n4063), .b(n3987), .O(n4077));
  orx  g4037(.a(n4077), .b(n4076), .O(n4078));
  andx g4038(.a(n4056), .b(n4003), .O(n4079));
  andx g4039(.a(n4021), .b(n3977), .O(n4080));
  orx  g4040(.a(n4080), .b(n4079), .O(n4081));
  orx  g4041(.a(n4081), .b(n4078), .O(n4082));
  orx  g4042(.a(n4082), .b(n4075), .O(n4083));
  orx  g4043(.a(n4083), .b(n4067), .O(n4084));
  orx  g4044(.a(n4084), .b(n4044), .O(n4085));
  orx  g4045(.a(n4085), .b(n3952), .O(n4086));
  andx g4046(.a(n3539), .b(n88), .O(n4087));
  andx g4047(.a(n43), .b(n3187), .O(n4088));
  andx g4048(.a(n4088), .b(n48), .O(n4089));
  andx g4049(.a(n4089), .b(n4087), .O(n4090));
  andx g4050(.a(n3989), .b(n4090), .O(n4091));
  andx g4051(.a(n3539), .b(n3187), .O(n4092));
  andx g4052(.a(n4092), .b(n2508), .O(n4093));
  andx g4053(.a(n4093), .b(n3989), .O(n4094));
  andx g4054(.a(n3543), .b(n313), .O(n4095));
  andx g4055(.a(n3986), .b(n3181), .O(n4096));
  andx g4056(.a(n4096), .b(n4095), .O(n4097));
  orx  g4057(.a(n4097), .b(n4094), .O(n4098));
  orx  g4058(.a(n4098), .b(n4091), .O(n4099));
  andx g4059(.a(n3663), .b(n533), .O(n4100));
  andx g4060(.a(n3181), .b(n303), .O(n4101));
  andx g4061(.a(n4101), .b(n3508), .O(n4102));
  andx g4062(.a(n4102), .b(n4100), .O(n4103));
  andx g4063(.a(n3609), .b(n64), .O(n4104));
  andx g4064(.a(n4104), .b(n88), .O(n4105));
  andx g4065(.a(n4105), .b(n3576), .O(n4106));
  orx  g4066(.a(n4106), .b(n4103), .O(n4107));
  andx g4067(.a(n3932), .b(pi18), .O(n4108));
  andx g4068(.a(n4108), .b(n3189), .O(n4109));
  andx g4069(.a(n3736), .b(n3180), .O(n4110));
  andx g4070(.a(n4110), .b(n3843), .O(n4111));
  andx g4071(.a(n4111), .b(n4109), .O(n4112));
  andx g4072(.a(n3225), .b(n1687), .O(n4113));
  andx g4073(.a(n92), .b(pi35), .O(n4114));
  andx g4074(.a(n4114), .b(n4113), .O(n4115));
  orx  g4075(.a(n4115), .b(n4112), .O(n4116));
  orx  g4076(.a(n4116), .b(n4107), .O(n4117));
  andx g4077(.a(n3489), .b(n533), .O(n4118));
  andx g4078(.a(n4118), .b(n3640), .O(n4119));
  andx g4079(.a(n47), .b(pi07), .O(n4120));
  andx g4080(.a(n4120), .b(n43), .O(n4121));
  andx g4081(.a(n4033), .b(n644), .O(n4122));
  andx g4082(.a(n4122), .b(n4121), .O(n4123));
  andx g4083(.a(n4123), .b(n3995), .O(n4124));
  andx g4084(.a(n4124), .b(n4017), .O(n4125));
  orx  g4085(.a(n4125), .b(n4119), .O(n4126));
  andx g4086(.a(n2507), .b(n46), .O(n4127));
  andx g4087(.a(n3255), .b(n73), .O(n4128));
  andx g4088(.a(n4128), .b(n4127), .O(n4129));
  andx g4089(.a(n4129), .b(n3981), .O(n4130));
  andx g4090(.a(n4130), .b(n4017), .O(n4131));
  andx g4091(.a(n3685), .b(pi18), .O(n4132));
  andx g4092(.a(n4132), .b(n3266), .O(n4133));
  andx g4093(.a(n3290), .b(n63), .O(n4134));
  andx g4094(.a(n3218), .b(n1768), .O(n4135));
  andx g4095(.a(n4135), .b(n4134), .O(n4136));
  andx g4096(.a(n4136), .b(n4133), .O(n4137));
  orx  g4097(.a(n4137), .b(n4131), .O(n4138));
  orx  g4098(.a(n4138), .b(n4126), .O(n4139));
  orx  g4099(.a(n4139), .b(n4117), .O(n4140));
  orx  g4100(.a(n4140), .b(n4099), .O(n4141));
  andx g4101(.a(n3319), .b(n41), .O(n4142));
  andx g4102(.a(n43), .b(pi19), .O(n4143));
  andx g4103(.a(n4143), .b(n48), .O(n4144));
  andx g4104(.a(n4144), .b(n4142), .O(n4145));
  andx g4105(.a(n4145), .b(n3989), .O(n4146));
  andx g4106(.a(n3540), .b(n3203), .O(n4147));
  andx g4107(.a(n4147), .b(n4087), .O(n4148));
  andx g4108(.a(n4148), .b(n4030), .O(n4149));
  orx  g4109(.a(n4149), .b(n4146), .O(n4150));
  andx g4110(.a(n3568), .b(pi35), .O(n4151));
  andx g4111(.a(n4151), .b(n3617), .O(n4152));
  andx g4112(.a(n4104), .b(n41), .O(n4153));
  andx g4113(.a(n3508), .b(n3203), .O(n4154));
  andx g4114(.a(n3420), .b(n303), .O(n4155));
  andx g4115(.a(n4155), .b(n4154), .O(n4156));
  andx g4116(.a(n4156), .b(n4153), .O(n4157));
  orx  g4117(.a(n4157), .b(n4152), .O(n4158));
  orx  g4118(.a(n4158), .b(n4150), .O(n4159));
  andx g4119(.a(n3214), .b(n895), .O(n4160));
  andx g4120(.a(n4160), .b(n378), .O(n4161));
  andx g4121(.a(n4161), .b(n4133), .O(n4162));
  andx g4122(.a(n3567), .b(n88), .O(n4163));
  andx g4123(.a(n3203), .b(n3188), .O(n4164));
  andx g4124(.a(n4164), .b(n4163), .O(n4165));
  andx g4125(.a(n4010), .b(n3385), .O(n4166));
  andx g4126(.a(n4166), .b(n4165), .O(n4167));
  orx  g4127(.a(n4167), .b(n4162), .O(n4168));
  andx g4128(.a(n3761), .b(n3719), .O(n4169));
  andx g4129(.a(n4169), .b(n3960), .O(n4170));
  andx g4130(.a(n303), .b(n75), .O(n4171));
  andx g4131(.a(n4171), .b(n3784), .O(n4172));
  andx g4132(.a(n4172), .b(n4170), .O(n4173));
  andx g4133(.a(n3732), .b(n3187), .O(n4174));
  andx g4134(.a(n3735), .b(n2544), .O(n4175));
  andx g4135(.a(n4175), .b(n4174), .O(n4176));
  andx g4136(.a(n4176), .b(n3250), .O(n4177));
  orx  g4137(.a(n4177), .b(n4173), .O(n4178));
  orx  g4138(.a(n4178), .b(n4168), .O(n4179));
  orx  g4139(.a(n4179), .b(n4159), .O(n4180));
  andx g4140(.a(n4123), .b(n4025), .O(n4181));
  andx g4141(.a(n4002), .b(n4181), .O(n4182));
  andx g4142(.a(n3187), .b(pi07), .O(n4183));
  andx g4143(.a(n4183), .b(n3735), .O(n4184));
  andx g4144(.a(n4184), .b(n3733), .O(n4185));
  andx g4145(.a(n4185), .b(n3471), .O(n4186));
  orx  g4146(.a(n4186), .b(n4182), .O(n4187));
  andx g4147(.a(n3319), .b(n88), .O(n4188));
  andx g4148(.a(n93), .b(pi19), .O(n4189));
  andx g4149(.a(n4189), .b(n3203), .O(n4190));
  andx g4150(.a(n4190), .b(n4188), .O(n4191));
  andx g4151(.a(n4191), .b(n3955), .O(n4192));
  andx g4152(.a(n3971), .b(n3255), .O(n4193));
  andx g4153(.a(n4193), .b(n4143), .O(n4194));
  andx g4154(.a(n4194), .b(n4163), .O(n4195));
  andx g4155(.a(n4195), .b(n3987), .O(n4196));
  orx  g4156(.a(n4196), .b(n4192), .O(n4197));
  orx  g4157(.a(n4197), .b(n4187), .O(n4198));
  andx g4158(.a(n3232), .b(n3193), .O(n4199));
  andx g4159(.a(n3290), .b(n3199), .O(n4200));
  andx g4160(.a(n4200), .b(n4199), .O(n4201));
  andx g4161(.a(n3567), .b(n3187), .O(n4202));
  andx g4162(.a(n41), .b(pi19), .O(n4203));
  andx g4163(.a(n4203), .b(n3203), .O(n4204));
  andx g4164(.a(n4204), .b(n4202), .O(n4205));
  andx g4165(.a(n4205), .b(n4201), .O(n4206));
  andx g4166(.a(n4190), .b(n4142), .O(n4207));
  andx g4167(.a(n4207), .b(n3955), .O(n4208));
  orx  g4168(.a(n4208), .b(n4206), .O(n4209));
  andx g4169(.a(n3270), .b(n3231), .O(n4210));
  andx g4170(.a(n4210), .b(n4113), .O(n4211));
  andx g4171(.a(n3469), .b(n91), .O(n4212));
  andx g4172(.a(n4212), .b(n3419), .O(n4213));
  andx g4173(.a(n4213), .b(n4100), .O(n4214));
  orx  g4174(.a(n4214), .b(n4211), .O(n4215));
  orx  g4175(.a(n4215), .b(n4209), .O(n4216));
  orx  g4176(.a(n4216), .b(n4198), .O(n4217));
  orx  g4177(.a(n4217), .b(n4180), .O(n4218));
  andx g4178(.a(n4169), .b(n3956), .O(n4219));
  andx g4179(.a(n4219), .b(n4172), .O(n4220));
  andx g4180(.a(n3871), .b(n3255), .O(n4221));
  andx g4181(.a(n4221), .b(n4143), .O(n4222));
  andx g4182(.a(n4222), .b(n4202), .O(n4223));
  andx g4183(.a(n4223), .b(n3987), .O(n4224));
  orx  g4184(.a(n4224), .b(n4220), .O(n4225));
  andx g4185(.a(n4176), .b(n3471), .O(n4226));
  andx g4186(.a(n3187), .b(n64), .O(n4227));
  andx g4187(.a(n4227), .b(n3203), .O(n4228));
  andx g4188(.a(n4228), .b(n3969), .O(n4229));
  andx g4189(.a(n4229), .b(n4201), .O(n4230));
  orx  g4190(.a(n4230), .b(n4226), .O(n4231));
  orx  g4191(.a(n4231), .b(n4225), .O(n4232));
  andx g4192(.a(n3736), .b(n313), .O(n4233));
  andx g4193(.a(n4233), .b(n3852), .O(n4234));
  andx g4194(.a(n4234), .b(n4109), .O(n4235));
  andx g4195(.a(n41), .b(n64), .O(n4236));
  andx g4196(.a(n4236), .b(n3203), .O(n4237));
  andx g4197(.a(n4237), .b(n3981), .O(n4238));
  andx g4198(.a(n4238), .b(n4201), .O(n4239));
  orx  g4199(.a(n4239), .b(n4235), .O(n4240));
  andx g4200(.a(n4132), .b(n3189), .O(n4241));
  andx g4201(.a(n3469), .b(n44), .O(n4242));
  andx g4202(.a(n3736), .b(n3181), .O(n4243));
  andx g4203(.a(n4243), .b(n4242), .O(n4244));
  andx g4204(.a(n4244), .b(n4241), .O(n4245));
  andx g4205(.a(n4153), .b(n3576), .O(n4246));
  orx  g4206(.a(n4246), .b(n4245), .O(n4247));
  orx  g4207(.a(n4247), .b(n4240), .O(n4248));
  orx  g4208(.a(n4248), .b(n4232), .O(n4249));
  andx g4209(.a(n4108), .b(n3266), .O(n4250));
  andx g4210(.a(n3374), .b(n3843), .O(n4251));
  andx g4211(.a(n4251), .b(n4250), .O(n4252));
  andx g4212(.a(n93), .b(n41), .O(n4253));
  andx g4213(.a(n4253), .b(n3203), .O(n4254));
  andx g4214(.a(n4254), .b(n4092), .O(n4255));
  andx g4215(.a(n4255), .b(n3955), .O(n4256));
  orx  g4216(.a(n4256), .b(n4252), .O(n4257));
  andx g4217(.a(n3784), .b(n1503), .O(n4258));
  andx g4218(.a(n4258), .b(n4095), .O(n4259));
  andx g4219(.a(n3288), .b(n644), .O(n4260));
  andx g4220(.a(n3698), .b(n3419), .O(n4261));
  andx g4221(.a(n4261), .b(n4260), .O(n4262));
  orx  g4222(.a(n4262), .b(n4259), .O(n4263));
  orx  g4223(.a(n4263), .b(n4257), .O(n4264));
  andx g4224(.a(n4238), .b(n4166), .O(n4265));
  andx g4225(.a(n4191), .b(n4030), .O(n4266));
  orx  g4226(.a(n4266), .b(n4265), .O(n4267));
  andx g4227(.a(n4151), .b(n3328), .O(n4268));
  andx g4228(.a(n3735), .b(n3203), .O(n4269));
  andx g4229(.a(n4269), .b(n3995), .O(n4270));
  andx g4230(.a(n4270), .b(n4201), .O(n4271));
  orx  g4231(.a(n4271), .b(n4268), .O(n4272));
  orx  g4232(.a(n4272), .b(n4267), .O(n4273));
  orx  g4233(.a(n4273), .b(n4264), .O(n4274));
  orx  g4234(.a(n4274), .b(n4249), .O(n4275));
  orx  g4235(.a(n4275), .b(n4218), .O(n4276));
  orx  g4236(.a(n4276), .b(n4141), .O(n4277));
  andx g4237(.a(n3566), .b(n3521), .O(n4278));
  andx g4238(.a(pi30), .b(pi12), .O(n4279));
  andx g4239(.a(n4279), .b(n200), .O(n4280));
  andx g4240(.a(n4280), .b(pi32), .O(n4281));
  orx  g4241(.a(n4281), .b(n4278), .O(n4282));
  andx g4242(.a(pi16), .b(n3193), .O(n4283));
  andx g4243(.a(n4283), .b(n3937), .O(n4284));
  andx g4244(.a(n4284), .b(n3321), .O(n4285));
  andx g4245(.a(n3290), .b(n644), .O(n4286));
  andx g4246(.a(n4286), .b(n4285), .O(n4287));
  andx g4247(.a(pi35), .b(pi09), .O(n4288));
  andx g4248(.a(n3427), .b(n42), .O(n4289));
  andx g4249(.a(n4289), .b(n4288), .O(n4290));
  andx g4250(.a(n3055), .b(n644), .O(n4291));
  andx g4251(.a(n4291), .b(n49), .O(n4292));
  andx g4252(.a(n4292), .b(n4290), .O(n4293));
  orx  g4253(.a(n4293), .b(n4287), .O(n4294));
  orx  g4254(.a(n4294), .b(n4282), .O(n4295));
  andx g4255(.a(pi20), .b(pi21), .O(n4296));
  andx g4256(.a(n4279), .b(n63), .O(n4297));
  andx g4257(.a(n4297), .b(n182), .O(n4298));
  andx g4258(.a(n4298), .b(n4296), .O(n4299));
  andx g4259(.a(pi16), .b(n87), .O(n4300));
  andx g4260(.a(n4300), .b(n1831), .O(n4301));
  andx g4261(.a(n4301), .b(n3321), .O(n4302));
  andx g4262(.a(n3818), .b(n4302), .O(n4303));
  orx  g4263(.a(n4303), .b(n4299), .O(n4304));
  andx g4264(.a(pi09), .b(pi29), .O(n4305));
  andx g4265(.a(n4305), .b(n333), .O(n4306));
  andx g4266(.a(n4306), .b(n437), .O(n4307));
  andx g4267(.a(n4307), .b(pi27), .O(n4308));
  andx g4268(.a(pi09), .b(pi12), .O(n4309));
  andx g4269(.a(n4309), .b(n1127), .O(n4310));
  andx g4270(.a(n4310), .b(n4296), .O(n4311));
  orx  g4271(.a(n4311), .b(n4308), .O(n4312));
  orx  g4272(.a(n4312), .b(n4304), .O(n4313));
  orx  g4273(.a(n4313), .b(n4295), .O(n4314));
  andx g4274(.a(n3188), .b(n449), .O(n4315));
  andx g4275(.a(n3305), .b(n431), .O(n4316));
  andx g4276(.a(n4316), .b(n4315), .O(n4317));
  andx g4277(.a(n4317), .b(n4102), .O(n4318));
  andx g4278(.a(n52), .b(n1687), .O(n4319));
  andx g4279(.a(n4319), .b(n3180), .O(n4320));
  andx g4280(.a(pi26), .b(n43), .O(n4321));
  andx g4281(.a(n4321), .b(n3241), .O(n4322));
  andx g4282(.a(n4322), .b(n4320), .O(n4323));
  andx g4283(.a(n1942), .b(n107), .O(n4324));
  andx g4284(.a(n4324), .b(n3667), .O(n4325));
  andx g4285(.a(n4325), .b(n4323), .O(n4326));
  orx  g4286(.a(n4326), .b(n4318), .O(n4327));
  andx g4287(.a(pi20), .b(n91), .O(n4328));
  andx g4288(.a(n4328), .b(n895), .O(n4329));
  andx g4289(.a(n4329), .b(n3271), .O(n4330));
  andx g4290(.a(n4330), .b(n3488), .O(n4331));
  orx  g4291(.a(n4331), .b(n384), .O(n4332));
  orx  g4292(.a(n4332), .b(n4327), .O(n4333));
  andx g4293(.a(n4288), .b(n63), .O(n4334));
  andx g4294(.a(n42), .b(n67), .O(n4335));
  andx g4295(.a(n4335), .b(n4334), .O(n4336));
  andx g4296(.a(n3367), .b(n2507), .O(n4337));
  andx g4297(.a(n3910), .b(n756), .O(n4338));
  andx g4298(.a(n4338), .b(n4337), .O(n4339));
  andx g4299(.a(n4339), .b(n4336), .O(n4340));
  andx g4300(.a(n855), .b(n75), .O(n4341));
  andx g4301(.a(n329), .b(n64), .O(n4342));
  andx g4302(.a(n4342), .b(n4341), .O(n4343));
  andx g4303(.a(n3508), .b(n3253), .O(n4344));
  andx g4304(.a(n3203), .b(n301), .O(n4345));
  andx g4305(.a(n4345), .b(n4344), .O(n4346));
  andx g4306(.a(n4346), .b(n4343), .O(n4347));
  orx  g4307(.a(n4347), .b(n4340), .O(n4348));
  andx g4308(.a(n3214), .b(n229), .O(n4349));
  andx g4309(.a(n533), .b(pi16), .O(n4350));
  andx g4310(.a(n4350), .b(n1901), .O(n4351));
  andx g4311(.a(n4351), .b(n4349), .O(n4352));
  andx g4312(.a(n4352), .b(n766), .O(n4353));
  andx g4313(.a(n64), .b(pi15), .O(n4354));
  andx g4314(.a(n4354), .b(pi16), .O(n4355));
  andx g4315(.a(n4355), .b(n3684), .O(n4356));
  andx g4316(.a(n3757), .b(n4356), .O(n4357));
  orx  g4317(.a(n4357), .b(n4353), .O(n4358));
  orx  g4318(.a(n4358), .b(n4348), .O(n4359));
  orx  g4319(.a(n4359), .b(n4333), .O(n4360));
  orx  g4320(.a(n4360), .b(n4314), .O(n4361));
  andx g4321(.a(n3855), .b(n855), .O(n4362));
  andx g4322(.a(n4362), .b(n1689), .O(n4363));
  andx g4323(.a(n4363), .b(n3344), .O(n4364));
  andx g4324(.a(n1815), .b(pi30), .O(n4365));
  andx g4325(.a(n4365), .b(n437), .O(n4366));
  andx g4326(.a(n4366), .b(n4296), .O(n4367));
  orx  g4327(.a(n4367), .b(n4364), .O(n4368));
  andx g4328(.a(n522), .b(n110), .O(n4369));
  andx g4329(.a(n4369), .b(pi32), .O(n4370));
  andx g4330(.a(n75), .b(pi08), .O(n4371));
  andx g4331(.a(n4371), .b(n522), .O(n4372));
  andx g4332(.a(n4372), .b(n4296), .O(n4373));
  orx  g4333(.a(n4373), .b(n4370), .O(n4374));
  orx  g4334(.a(n4374), .b(n4368), .O(n4375));
  andx g4335(.a(n4057), .b(n285), .O(n4376));
  andx g4336(.a(n4376), .b(pi27), .O(n4377));
  andx g4337(.a(n4296), .b(n4280), .O(n4378));
  orx  g4338(.a(n4378), .b(n4377), .O(n4379));
  andx g4339(.a(n4302), .b(n4160), .O(n4380));
  andx g4340(.a(n75), .b(pi12), .O(n4381));
  andx g4341(.a(n4381), .b(n522), .O(n4382));
  andx g4342(.a(n4382), .b(pi32), .O(n4383));
  orx  g4343(.a(n4383), .b(n4380), .O(n4384));
  orx  g4344(.a(n4384), .b(n4379), .O(n4385));
  orx  g4345(.a(n4385), .b(n4375), .O(n4386));
  andx g4346(.a(n4376), .b(pi28), .O(n4387));
  andx g4347(.a(pi09), .b(pi08), .O(n4388));
  andx g4348(.a(n4388), .b(n1127), .O(n4389));
  andx g4349(.a(n4389), .b(n4296), .O(n4390));
  orx  g4350(.a(n4390), .b(n4387), .O(n4391));
  andx g4351(.a(n3856), .b(n3290), .O(n4392));
  andx g4352(.a(n4392), .b(n3843), .O(n4393));
  andx g4353(.a(n4393), .b(n3391), .O(n4394));
  andx g4354(.a(pi30), .b(pi08), .O(n4395));
  andx g4355(.a(n4395), .b(n200), .O(n4396));
  andx g4356(.a(n4396), .b(pi32), .O(n4397));
  orx  g4357(.a(n4397), .b(n4394), .O(n4398));
  orx  g4358(.a(n4398), .b(n4391), .O(n4399));
  andx g4359(.a(n3270), .b(n91), .O(n4400));
  andx g4360(.a(n3462), .b(n3419), .O(n4401));
  andx g4361(.a(n4401), .b(n4400), .O(n4402));
  andx g4362(.a(n4402), .b(n3662), .O(n4403));
  andx g4363(.a(n3469), .b(n430), .O(n4404));
  andx g4364(.a(n4404), .b(n4285), .O(n4405));
  orx  g4365(.a(n4405), .b(n4403), .O(n4406));
  andx g4366(.a(pi11), .b(n63), .O(n4407));
  andx g4367(.a(n4407), .b(pi30), .O(n4408));
  andx g4368(.a(n4408), .b(n182), .O(n4409));
  andx g4369(.a(n4409), .b(n4296), .O(n4410));
  andx g4370(.a(n3855), .b(n1689), .O(n4411));
  andx g4371(.a(n4411), .b(n3419), .O(n4412));
  andx g4372(.a(n4412), .b(n3224), .O(n4413));
  orx  g4373(.a(n4413), .b(n4410), .O(n4414));
  orx  g4374(.a(n4414), .b(n4406), .O(n4415));
  orx  g4375(.a(n4415), .b(n4399), .O(n4416));
  orx  g4376(.a(n4416), .b(n4386), .O(n4417));
  orx  g4377(.a(n4417), .b(n4361), .O(n4418));
  andx g4378(.a(n4350), .b(n64), .O(n4419));
  andx g4379(.a(n4419), .b(n3608), .O(n4420));
  andx g4380(.a(n3806), .b(n4420), .O(n4421));
  orx  g4381(.a(n4421), .b(n1864), .O(n4422));
  andx g4382(.a(n3180), .b(n756), .O(n4423));
  andx g4383(.a(n3382), .b(n3259), .O(n4424));
  andx g4384(.a(n4424), .b(n4423), .O(n4425));
  andx g4385(.a(n3556), .b(n3367), .O(n4426));
  andx g4386(.a(n4426), .b(n4324), .O(n4427));
  andx g4387(.a(n4427), .b(n4425), .O(n4428));
  andx g4388(.a(n2682), .b(n313), .O(n4429));
  andx g4389(.a(n4429), .b(n2909), .O(n4430));
  andx g4390(.a(n199), .b(n107), .O(n4431));
  andx g4391(.a(n4431), .b(n3734), .O(n4432));
  andx g4392(.a(n4432), .b(n4430), .O(n4433));
  orx  g4393(.a(n4433), .b(n4428), .O(n4434));
  orx  g4394(.a(n4434), .b(n4422), .O(n4435));
  andx g4395(.a(n229), .b(n42), .O(n4436));
  andx g4396(.a(n4436), .b(n3469), .O(n4437));
  andx g4397(.a(n73), .b(n45), .O(n4438));
  andx g4398(.a(n4438), .b(n3602), .O(n4439));
  andx g4399(.a(n4439), .b(n4437), .O(n4440));
  andx g4400(.a(n3428), .b(n229), .O(n4441));
  andx g4401(.a(n4441), .b(n3290), .O(n4442));
  andx g4402(.a(n47), .b(n249), .O(n4443));
  andx g4403(.a(n4443), .b(n3253), .O(n4444));
  andx g4404(.a(n2507), .b(n644), .O(n4445));
  andx g4405(.a(n4445), .b(n4444), .O(n4446));
  andx g4406(.a(n4446), .b(n4442), .O(n4447));
  orx  g4407(.a(n4447), .b(n4440), .O(n4448));
  andx g4408(.a(n3772), .b(n3218), .O(n4449));
  andx g4409(.a(n4449), .b(n3480), .O(n4450));
  andx g4410(.a(n4450), .b(n3662), .O(n4451));
  andx g4411(.a(n3305), .b(n3239), .O(n4452));
  andx g4412(.a(n4452), .b(n4315), .O(n4453));
  andx g4413(.a(n3699), .b(n4453), .O(n4454));
  orx  g4414(.a(n4454), .b(n4451), .O(n4455));
  orx  g4415(.a(n4455), .b(n4448), .O(n4456));
  orx  g4416(.a(n4456), .b(n4435), .O(n4457));
  andx g4417(.a(n4441), .b(n895), .O(n4458));
  andx g4418(.a(n3719), .b(n48), .O(n4459));
  andx g4419(.a(n4459), .b(n3220), .O(n4460));
  andx g4420(.a(n4460), .b(n4458), .O(n4461));
  andx g4421(.a(n644), .b(n437), .O(n4462));
  andx g4422(.a(n4462), .b(n4288), .O(n4463));
  andx g4423(.a(n107), .b(n1687), .O(n4464));
  andx g4424(.a(n4464), .b(n45), .O(n4465));
  andx g4425(.a(n533), .b(n42), .O(n4466));
  andx g4426(.a(n4466), .b(n48), .O(n4467));
  andx g4427(.a(n4467), .b(n4465), .O(n4468));
  andx g4428(.a(n4468), .b(n4463), .O(n4469));
  orx  g4429(.a(n4469), .b(n4461), .O(n4470));
  andx g4430(.a(n3214), .b(n357), .O(n4471));
  andx g4431(.a(n4471), .b(n2508), .O(n4472));
  andx g4432(.a(n4472), .b(n4458), .O(n4473));
  andx g4433(.a(n3621), .b(n3331), .O(n4474));
  orx  g4434(.a(n4474), .b(n4473), .O(n4475));
  orx  g4435(.a(n4475), .b(n4470), .O(n4476));
  andx g4436(.a(n4289), .b(n381), .O(n4477));
  andx g4437(.a(n3624), .b(n48), .O(n4478));
  andx g4438(.a(n756), .b(n45), .O(n4479));
  andx g4439(.a(n4479), .b(n4478), .O(n4480));
  andx g4440(.a(n4480), .b(n4477), .O(n4481));
  andx g4441(.a(n3219), .b(n48), .O(n4482));
  andx g4442(.a(n4482), .b(n4479), .O(n4483));
  andx g4443(.a(n4483), .b(n4477), .O(n4484));
  orx  g4444(.a(n4484), .b(n4481), .O(n4485));
  andx g4445(.a(n3695), .b(n1344), .O(n4486));
  andx g4446(.a(n1768), .b(n1688), .O(n4487));
  andx g4447(.a(n4487), .b(n4134), .O(n4488));
  andx g4448(.a(n4488), .b(n4486), .O(n4489));
  orx  g4449(.a(n4489), .b(n1533), .O(n4490));
  orx  g4450(.a(n4490), .b(n4485), .O(n4491));
  orx  g4451(.a(n4491), .b(n4476), .O(n4492));
  orx  g4452(.a(n4492), .b(n4457), .O(n4493));
  andx g4453(.a(n3403), .b(pi07), .O(n4494));
  andx g4454(.a(n4494), .b(n4341), .O(n4495));
  andx g4455(.a(n345), .b(n298), .O(n4496));
  andx g4456(.a(n4443), .b(n3246), .O(n4497));
  andx g4457(.a(n4497), .b(n4496), .O(n4498));
  andx g4458(.a(n4498), .b(n4495), .O(n4499));
  andx g4459(.a(n3241), .b(n313), .O(n4500));
  andx g4460(.a(n4319), .b(n2256), .O(n4501));
  andx g4461(.a(n4501), .b(n4500), .O(n4502));
  andx g4462(.a(n4502), .b(n4432), .O(n4503));
  orx  g4463(.a(n4503), .b(n4499), .O(n4504));
  andx g4464(.a(n4497), .b(n4445), .O(n4505));
  andx g4465(.a(n4505), .b(n4495), .O(n4506));
  andx g4466(.a(n3566), .b(n3331), .O(n4507));
  orx  g4467(.a(n4507), .b(n4506), .O(n4508));
  orx  g4468(.a(n4508), .b(n4504), .O(n4509));
  andx g4469(.a(n3314), .b(n756), .O(n4510));
  andx g4470(.a(n4510), .b(n3552), .O(n4511));
  andx g4471(.a(n4511), .b(n3558), .O(n4512));
  andx g4472(.a(n3621), .b(n3521), .O(n4513));
  orx  g4473(.a(n4513), .b(n4512), .O(n4514));
  andx g4474(.a(n2964), .b(n229), .O(n4515));
  andx g4475(.a(n4350), .b(n644), .O(n4516));
  andx g4476(.a(n4516), .b(n4515), .O(n4517));
  andx g4477(.a(n4517), .b(n3480), .O(n4518));
  andx g4478(.a(n3688), .b(n4356), .O(n4519));
  orx  g4479(.a(n4519), .b(n4518), .O(n4520));
  orx  g4480(.a(n4520), .b(n4514), .O(n4521));
  orx  g4481(.a(n4521), .b(n4509), .O(n4522));
  andx g4482(.a(n4354), .b(n3644), .O(n4523));
  andx g4483(.a(n3305), .b(n229), .O(n4524));
  andx g4484(.a(n4524), .b(n4523), .O(n4525));
  andx g4485(.a(n4525), .b(n4102), .O(n4526));
  orx  g4486(.a(n4526), .b(n1715), .O(n4527));
  andx g4487(.a(n4511), .b(n3668), .O(n4528));
  andx g4488(.a(n4496), .b(n4444), .O(n4529));
  andx g4489(.a(n4529), .b(n4442), .O(n4530));
  orx  g4490(.a(n4530), .b(n4528), .O(n4531));
  orx  g4491(.a(n4531), .b(n4527), .O(n4532));
  andx g4492(.a(n4213), .b(n4317), .O(n4533));
  andx g4493(.a(n4321), .b(n4319), .O(n4534));
  andx g4494(.a(n4534), .b(n4500), .O(n4535));
  andx g4495(.a(n4431), .b(n3605), .O(n4536));
  andx g4496(.a(n4536), .b(n4535), .O(n4537));
  orx  g4497(.a(n4537), .b(n4533), .O(n4538));
  andx g4498(.a(n4328), .b(n1021), .O(n4539));
  andx g4499(.a(n4539), .b(n4134), .O(n4540));
  andx g4500(.a(n4540), .b(n3488), .O(n4541));
  andx g4501(.a(n3234), .b(n75), .O(n4542));
  andx g4502(.a(n4542), .b(n3403), .O(n4543));
  andx g4503(.a(n2544), .b(n644), .O(n4544));
  andx g4504(.a(n4544), .b(n49), .O(n4545));
  andx g4505(.a(n4545), .b(n4543), .O(n4546));
  orx  g4506(.a(n4546), .b(n4541), .O(n4547));
  orx  g4507(.a(n4547), .b(n4538), .O(n4548));
  orx  g4508(.a(n4548), .b(n4532), .O(n4549));
  orx  g4509(.a(n4549), .b(n4522), .O(n4550));
  orx  g4510(.a(n4550), .b(n4493), .O(n4551));
  orx  g4511(.a(n4551), .b(n4418), .O(n4552));
  andx g4512(.a(n4396), .b(n4296), .O(n4553));
  andx g4513(.a(n4280), .b(pi33), .O(n4554));
  orx  g4514(.a(n4554), .b(n4553), .O(n4555));
  andx g4515(.a(n4307), .b(pi28), .O(n4556));
  andx g4516(.a(n4396), .b(pi33), .O(n4557));
  orx  g4517(.a(n4557), .b(n4556), .O(n4558));
  orx  g4518(.a(n4558), .b(n4555), .O(n4559));
  andx g4519(.a(n4366), .b(pi33), .O(n4560));
  andx g4520(.a(n313), .b(n1687), .O(n4561));
  andx g4521(.a(n1344), .b(n65), .O(n4562));
  andx g4522(.a(n4562), .b(n3855), .O(n4563));
  andx g4523(.a(n4563), .b(n4561), .O(n4564));
  orx  g4524(.a(n4564), .b(n4560), .O(n4565));
  andx g4525(.a(n3224), .b(n3183), .O(n4566));
  andx g4526(.a(n3427), .b(n75), .O(n4567));
  andx g4527(.a(n4567), .b(n1901), .O(n4568));
  andx g4528(.a(n3180), .b(n73), .O(n4569));
  andx g4529(.a(n4569), .b(n4568), .O(n4570));
  orx  g4530(.a(n4570), .b(n4566), .O(n4571));
  orx  g4531(.a(n4571), .b(n4565), .O(n4572));
  orx  g4532(.a(n4572), .b(n4559), .O(n4573));
  andx g4533(.a(n1815), .b(n1127), .O(n4574));
  andx g4534(.a(n4574), .b(pi33), .O(n4575));
  andx g4535(.a(n4382), .b(pi33), .O(n4576));
  orx  g4536(.a(n4576), .b(n4575), .O(n4577));
  andx g4537(.a(n4366), .b(pi32), .O(n4578));
  andx g4538(.a(n1081), .b(n333), .O(n4579));
  andx g4539(.a(n4579), .b(pi32), .O(n4580));
  orx  g4540(.a(n4580), .b(n4578), .O(n4581));
  orx  g4541(.a(n4581), .b(n4577), .O(n4582));
  andx g4542(.a(n4369), .b(pi33), .O(n4583));
  orx  g4543(.a(n4583), .b(n1434), .O(n4584));
  andx g4544(.a(n4389), .b(pi32), .O(n4585));
  orx  g4545(.a(n4585), .b(n2088), .O(n4586));
  orx  g4546(.a(n4586), .b(n4584), .O(n4587));
  orx  g4547(.a(n4587), .b(n4582), .O(n4588));
  orx  g4548(.a(n4588), .b(n4573), .O(n4589));
  andx g4549(.a(n756), .b(n484), .O(n4590));
  andx g4550(.a(n4590), .b(n49), .O(n4591));
  andx g4551(.a(n4591), .b(n4290), .O(n4592));
  andx g4552(.a(n3422), .b(n3253), .O(n4593));
  andx g4553(.a(n345), .b(n45), .O(n4594));
  andx g4554(.a(n4594), .b(n4593), .O(n4595));
  andx g4555(.a(n4595), .b(n3526), .O(n4596));
  orx  g4556(.a(n4596), .b(n4592), .O(n4597));
  andx g4557(.a(n230), .b(n1901), .O(n4598));
  andx g4558(.a(n3419), .b(pi35), .O(n4599));
  andx g4559(.a(n4599), .b(n357), .O(n4600));
  andx g4560(.a(n4600), .b(n4598), .O(n4601));
  andx g4561(.a(n3821), .b(n92), .O(n4602));
  andx g4562(.a(n4602), .b(n756), .O(n4603));
  andx g4563(.a(n4603), .b(n1966), .O(n4604));
  orx  g4564(.a(n4604), .b(n4601), .O(n4605));
  orx  g4565(.a(n4605), .b(n4597), .O(n4606));
  andx g4566(.a(n3193), .b(n91), .O(n4607));
  andx g4567(.a(n44), .b(n52), .O(n4608));
  andx g4568(.a(n4608), .b(n4607), .O(n4609));
  andx g4569(.a(n4609), .b(n644), .O(n4610));
  andx g4570(.a(n4610), .b(n4334), .O(n4611));
  orx  g4571(.a(n4611), .b(n340), .O(n4612));
  andx g4572(.a(n44), .b(pi07), .O(n4613));
  andx g4573(.a(n4613), .b(n1768), .O(n4614));
  andx g4574(.a(n4614), .b(n449), .O(n4615));
  andx g4575(.a(n4615), .b(n3687), .O(n4616));
  andx g4576(.a(n42), .b(pi09), .O(n4617));
  andx g4577(.a(n4617), .b(n3687), .O(n4618));
  andx g4578(.a(n4618), .b(n4591), .O(n4619));
  orx  g4579(.a(n4619), .b(n4616), .O(n4620));
  orx  g4580(.a(n4620), .b(n4612), .O(n4621));
  orx  g4581(.a(n4621), .b(n4606), .O(n4622));
  andx g4582(.a(n4389), .b(pi33), .O(n4623));
  andx g4583(.a(n3194), .b(n313), .O(n4624));
  andx g4584(.a(n4624), .b(n3855), .O(n4625));
  andx g4585(.a(n4625), .b(n522), .O(n4626));
  orx  g4586(.a(n4626), .b(n4623), .O(n4627));
  andx g4587(.a(n4369), .b(n4296), .O(n4628));
  andx g4588(.a(pi08), .b(n63), .O(n4629));
  andx g4589(.a(n4629), .b(pi30), .O(n4630));
  andx g4590(.a(n4630), .b(n182), .O(n4631));
  andx g4591(.a(n4631), .b(pi33), .O(n4632));
  orx  g4592(.a(n4632), .b(n4628), .O(n4633));
  orx  g4593(.a(n4633), .b(n4627), .O(n4634));
  andx g4594(.a(n73), .b(n1687), .O(n4635));
  andx g4595(.a(n3545), .b(n229), .O(n4636));
  andx g4596(.a(n4636), .b(n4635), .O(n4637));
  andx g4597(.a(n1773), .b(n756), .O(n4638));
  andx g4598(.a(n4638), .b(n49), .O(n4639));
  andx g4599(.a(n4639), .b(n4336), .O(n4640));
  orx  g4600(.a(n4640), .b(n4637), .O(n4641));
  andx g4601(.a(n4310), .b(pi33), .O(n4642));
  andx g4602(.a(n4579), .b(pi33), .O(n4643));
  orx  g4603(.a(n4643), .b(n4642), .O(n4644));
  orx  g4604(.a(n4644), .b(n4641), .O(n4645));
  orx  g4605(.a(n4645), .b(n4634), .O(n4646));
  orx  g4606(.a(n4646), .b(n4622), .O(n4647));
  orx  g4607(.a(n4647), .b(n4589), .O(n4648));
  andx g4608(.a(n4409), .b(pi32), .O(n4649));
  orx  g4609(.a(n4649), .b(n1419), .O(n4650));
  andx g4610(.a(n4183), .b(n538), .O(n4651));
  andx g4611(.a(n3786), .b(n229), .O(n4652));
  andx g4612(.a(n4652), .b(n4651), .O(n4653));
  andx g4613(.a(n4213), .b(n4653), .O(n4654));
  andx g4614(.a(n3843), .b(n3291), .O(n4655));
  andx g4615(.a(n4655), .b(n3696), .O(n4656));
  orx  g4616(.a(n4656), .b(n4654), .O(n4657));
  orx  g4617(.a(n4657), .b(n4650), .O(n4658));
  andx g4618(.a(n4213), .b(n4525), .O(n4659));
  andx g4619(.a(n4618), .b(n4292), .O(n4660));
  orx  g4620(.a(n4660), .b(n4659), .O(n4661));
  andx g4621(.a(n3180), .b(n1688), .O(n4662));
  andx g4622(.a(n4662), .b(n4598), .O(n4663));
  andx g4623(.a(n3910), .b(n73), .O(n4664));
  andx g4624(.a(n4664), .b(n3625), .O(n4665));
  andx g4625(.a(n4665), .b(n3404), .O(n4666));
  orx  g4626(.a(n4666), .b(n4663), .O(n4667));
  orx  g4627(.a(n4667), .b(n4661), .O(n4668));
  orx  g4628(.a(n4668), .b(n4658), .O(n4669));
  andx g4629(.a(n1688), .b(n1021), .O(n4670));
  andx g4630(.a(n1706), .b(n1454), .O(n4671));
  andx g4631(.a(n4671), .b(n3290), .O(n4672));
  andx g4632(.a(n4672), .b(n4670), .O(n4673));
  andx g4633(.a(n3856), .b(n895), .O(n4674));
  andx g4634(.a(n4674), .b(n3215), .O(n4675));
  andx g4635(.a(n4675), .b(n3706), .O(n4676));
  orx  g4636(.a(n4676), .b(n4673), .O(n4677));
  andx g4637(.a(n4382), .b(n4296), .O(n4678));
  andx g4638(.a(n4420), .b(n3516), .O(n4679));
  orx  g4639(.a(n4679), .b(n4678), .O(n4680));
  orx  g4640(.a(n4680), .b(n4677), .O(n4681));
  andx g4641(.a(n3321), .b(n3239), .O(n4682));
  andx g4642(.a(n3180), .b(n644), .O(n4683));
  andx g4643(.a(n4683), .b(n4682), .O(n4684));
  andx g4644(.a(n4542), .b(n329), .O(n4685));
  andx g4645(.a(n3881), .b(n48), .O(n4686));
  andx g4646(.a(n4236), .b(n313), .O(n4687));
  andx g4647(.a(n4687), .b(n4686), .O(n4688));
  andx g4648(.a(n4688), .b(n4685), .O(n4689));
  orx  g4649(.a(n4689), .b(n4684), .O(n4690));
  andx g4650(.a(n4372), .b(pi32), .O(n4691));
  orx  g4651(.a(n4691), .b(n2098), .O(n4692));
  orx  g4652(.a(n4692), .b(n4690), .O(n4693));
  orx  g4653(.a(n4693), .b(n4681), .O(n4694));
  orx  g4654(.a(n4694), .b(n4669), .O(n4695));
  andx g4655(.a(n4574), .b(pi32), .O(n4696));
  andx g4656(.a(n4631), .b(pi32), .O(n4697));
  orx  g4657(.a(n4697), .b(n4696), .O(n4698));
  andx g4658(.a(n4653), .b(n4102), .O(n4699));
  andx g4659(.a(n4409), .b(pi33), .O(n4700));
  orx  g4660(.a(n4700), .b(n4699), .O(n4701));
  orx  g4661(.a(n4701), .b(n4698), .O(n4702));
  andx g4662(.a(n3342), .b(n4486), .O(n4703));
  andx g4663(.a(n4372), .b(pi33), .O(n4704));
  orx  g4664(.a(n4704), .b(n4703), .O(n4705));
  andx g4665(.a(n4631), .b(n4296), .O(n4706));
  andx g4666(.a(n4574), .b(n4296), .O(n4707));
  orx  g4667(.a(n4707), .b(n4706), .O(n4708));
  orx  g4668(.a(n4708), .b(n4705), .O(n4709));
  orx  g4669(.a(n4709), .b(n4702), .O(n4710));
  andx g4670(.a(n4298), .b(pi32), .O(n4711));
  andx g4671(.a(n4579), .b(n4296), .O(n4712));
  orx  g4672(.a(n4712), .b(n4711), .O(n4713));
  andx g4673(.a(n4298), .b(pi33), .O(n4714));
  andx g4674(.a(n4310), .b(pi32), .O(n4715));
  orx  g4675(.a(n4715), .b(n4714), .O(n4716));
  orx  g4676(.a(n4716), .b(n4713), .O(n4717));
  andx g4677(.a(n3910), .b(n1688), .O(n4718));
  andx g4678(.a(n4718), .b(n3625), .O(n4719));
  andx g4679(.a(n4719), .b(n3526), .O(n4720));
  andx g4680(.a(n3246), .b(n3218), .O(n4721));
  andx g4681(.a(n3203), .b(n484), .O(n4722));
  andx g4682(.a(n4722), .b(n4721), .O(n4723));
  andx g4683(.a(n4723), .b(n4343), .O(n4724));
  orx  g4684(.a(n4724), .b(n4720), .O(n4725));
  andx g4685(.a(n3180), .b(n164), .O(n4726));
  andx g4686(.a(n4726), .b(n4682), .O(n4727));
  andx g4687(.a(n3508), .b(n65), .O(n4728));
  andx g4688(.a(n4728), .b(n3465), .O(n4729));
  andx g4689(.a(n4729), .b(n3696), .O(n4730));
  orx  g4690(.a(n4730), .b(n4727), .O(n4731));
  orx  g4691(.a(n4731), .b(n4725), .O(n4732));
  orx  g4692(.a(n4732), .b(n4717), .O(n4733));
  orx  g4693(.a(n4733), .b(n4710), .O(n4734));
  orx  g4694(.a(n4734), .b(n4695), .O(n4735));
  orx  g4695(.a(n4735), .b(n4648), .O(n4736));
  orx  g4696(.a(n4736), .b(n4552), .O(n4737));
  andx g4697(.a(n4201), .b(n4165), .O(n4738));
  andx g4698(.a(n3540), .b(n73), .O(n4739));
  andx g4699(.a(n4739), .b(n922), .O(n4740));
  andx g4700(.a(n4740), .b(n3969), .O(n4741));
  andx g4701(.a(n4741), .b(n4002), .O(n4742));
  orx  g4702(.a(n4742), .b(n4738), .O(n4743));
  andx g4703(.a(n4145), .b(n4039), .O(n4744));
  andx g4704(.a(n4205), .b(n4166), .O(n4745));
  orx  g4705(.a(n4745), .b(n4744), .O(n4746));
  orx  g4706(.a(n4746), .b(n4743), .O(n4747));
  andx g4707(.a(n1942), .b(n87), .O(n4748));
  andx g4708(.a(n4166), .b(n4270), .O(n4749));
  andx g4709(.a(n4188), .b(n4144), .O(n4750));
  andx g4710(.a(n4750), .b(n4039), .O(n4751));
  orx  g4711(.a(n4751), .b(n4749), .O(n4752));
  andx g4712(.a(n3861), .b(pi35), .O(n4753));
  andx g4713(.a(n4753), .b(n3328), .O(n4754));
  andx g4714(.a(n4181), .b(n4017), .O(n4755));
  orx  g4715(.a(n4755), .b(n4754), .O(n4756));
  orx  g4716(.a(n4756), .b(n4752), .O(n4757));
  orx  g4717(.a(n4757), .b(n4747), .O(n4758));
  andx g4718(.a(n4090), .b(n4039), .O(n4759));
  andx g4719(.a(n4156), .b(n4105), .O(n4760));
  orx  g4720(.a(n4760), .b(n4759), .O(n4761));
  andx g4721(.a(n3821), .b(n3340), .O(n4762));
  andx g4722(.a(n4762), .b(n4260), .O(n4763));
  andx g4723(.a(n4753), .b(n3617), .O(n4764));
  orx  g4724(.a(n4764), .b(n4763), .O(n4765));
  orx  g4725(.a(n4765), .b(n4761), .O(n4766));
  andx g4726(.a(n3270), .b(n1768), .O(n4767));
  andx g4727(.a(n4767), .b(n3393), .O(n4768));
  andx g4728(.a(n4768), .b(n4250), .O(n4769));
  andx g4729(.a(n4185), .b(n3250), .O(n4770));
  orx  g4730(.a(n4770), .b(n4769), .O(n4771));
  andx g4731(.a(n4233), .b(n3215), .O(n4772));
  andx g4732(.a(n4772), .b(n4241), .O(n4773));
  andx g4733(.a(n4229), .b(n4166), .O(n4774));
  orx  g4734(.a(n4774), .b(n4773), .O(n4775));
  orx  g4735(.a(n4775), .b(n4771), .O(n4776));
  orx  g4736(.a(n4776), .b(n4766), .O(n4777));
  orx  g4737(.a(n4777), .b(n4758), .O(n4778));
  andx g4738(.a(n4207), .b(n4030), .O(n4779));
  andx g4739(.a(n4002), .b(n4130), .O(n4780));
  orx  g4740(.a(n4780), .b(n4779), .O(n4781));
  andx g4741(.a(n4255), .b(n4030), .O(n4782));
  andx g4742(.a(n4002), .b(n4124), .O(n4783));
  orx  g4743(.a(n4783), .b(n4782), .O(n4784));
  orx  g4744(.a(n4784), .b(n4781), .O(n4785));
  andx g4745(.a(n4741), .b(n4017), .O(n4786));
  andx g4746(.a(n4453), .b(n3640), .O(n4787));
  andx g4747(.a(n4436), .b(n3214), .O(n4788));
  andx g4748(.a(n4545), .b(n4788), .O(n4789));
  orx  g4749(.a(n4789), .b(n4787), .O(n4790));
  orx  g4750(.a(n4790), .b(n1401), .O(n4791));
  orx  g4751(.a(n4791), .b(n4786), .O(n4792));
  andx g4752(.a(n4269), .b(n4025), .O(n4793));
  andx g4753(.a(n4793), .b(n4201), .O(n4794));
  andx g4754(.a(n4542), .b(n3419), .O(n4795));
  andx g4755(.a(n4795), .b(n4219), .O(n4796));
  orx  g4756(.a(n4796), .b(n4794), .O(n4797));
  orx  g4757(.a(n4797), .b(n4792), .O(n4798));
  orx  g4758(.a(n4798), .b(n4785), .O(n4799));
  andx g4759(.a(n4093), .b(n4039), .O(n4800));
  andx g4760(.a(n4793), .b(n4166), .O(n4801));
  orx  g4761(.a(n4801), .b(n4800), .O(n4802));
  andx g4762(.a(n3955), .b(n4148), .O(n4803));
  andx g4763(.a(n4223), .b(n4014), .O(n4804));
  orx  g4764(.a(n4804), .b(n4803), .O(n4805));
  orx  g4765(.a(n4805), .b(n4802), .O(n4806));
  andx g4766(.a(n4195), .b(n4014), .O(n4807));
  andx g4767(.a(n4118), .b(n3699), .O(n4808));
  orx  g4768(.a(n4808), .b(n4807), .O(n4809));
  andx g4769(.a(n4795), .b(n4170), .O(n4810));
  andx g4770(.a(n4750), .b(n3989), .O(n4811));
  orx  g4771(.a(n4811), .b(n4810), .O(n4812));
  orx  g4772(.a(n4812), .b(n4809), .O(n4813));
  orx  g4773(.a(n4813), .b(n4806), .O(n4814));
  orx  g4774(.a(n4814), .b(n4799), .O(n4815));
  orx  g4775(.a(n4815), .b(n4778), .O(n4816));
  orx  g4776(.a(n4816), .b(n4737), .O(n4817));
  andx g4777(.a(n4189), .b(n3319), .O(n4818));
  andx g4778(.a(n4818), .b(n3537), .O(n4819));
  andx g4779(.a(n3731), .b(n3705), .O(n4820));
  andx g4780(.a(n4820), .b(n3187), .O(n4821));
  andx g4781(.a(n3735), .b(n3255), .O(n4822));
  andx g4782(.a(n3406), .b(n2507), .O(n4823));
  andx g4783(.a(n4823), .b(n4822), .O(n4824));
  andx g4784(.a(n4824), .b(n3687), .O(n4825));
  andx g4785(.a(n4825), .b(n4821), .O(n4826));
  orx  g4786(.a(n4826), .b(n4819), .O(n4827));
  andx g4787(.a(n4324), .b(n3577), .O(n4828));
  andx g4788(.a(n3937), .b(n3422), .O(n4829));
  andx g4789(.a(n4829), .b(n3719), .O(n4830));
  andx g4790(.a(n4830), .b(n3421), .O(n4831));
  andx g4791(.a(n4831), .b(n4828), .O(n4832));
  andx g4792(.a(n3898), .b(n3234), .O(n4833));
  andx g4793(.a(n4443), .b(n3719), .O(n4834));
  andx g4794(.a(n4834), .b(n4833), .O(n4835));
  andx g4795(.a(n4835), .b(n3385), .O(n4836));
  andx g4796(.a(n4836), .b(n3197), .O(n4837));
  orx  g4797(.a(n4837), .b(n4832), .O(n4838));
  orx  g4798(.a(n4838), .b(n4827), .O(n4839));
  andx g4799(.a(n3855), .b(n3239), .O(n4840));
  andx g4800(.a(n4840), .b(n895), .O(n4841));
  andx g4801(.a(n4841), .b(n4057), .O(n4842));
  andx g4802(.a(n4842), .b(n3788), .O(n4843));
  andx g4803(.a(n3910), .b(pi35), .O(n4844));
  andx g4804(.a(n3882), .b(n73), .O(n4845));
  andx g4805(.a(n4845), .b(n4844), .O(n4846));
  andx g4806(.a(n4846), .b(n4828), .O(n4847));
  orx  g4807(.a(n4847), .b(n4843), .O(n4848));
  andx g4808(.a(n3872), .b(n3527), .O(n4849));
  andx g4809(.a(n3821), .b(n3231), .O(n4850));
  andx g4810(.a(n4850), .b(n230), .O(n4851));
  andx g4811(.a(n4851), .b(n3541), .O(n4852));
  orx  g4812(.a(n4852), .b(n4849), .O(n4853));
  orx  g4813(.a(n4853), .b(n4848), .O(n4854));
  orx  g4814(.a(n4854), .b(n4839), .O(n4855));
  andx g4815(.a(n3446), .b(n3334), .O(n4856));
  andx g4816(.a(n3609), .b(n88), .O(n4857));
  andx g4817(.a(n4857), .b(n3607), .O(n4858));
  orx  g4818(.a(n4858), .b(n4856), .O(n4859));
  andx g4819(.a(n3697), .b(n3640), .O(n4860));
  andx g4820(.a(n4682), .b(n64), .O(n4861));
  andx g4821(.a(n3290), .b(n1021), .O(n4862));
  andx g4822(.a(n4862), .b(n4861), .O(n4863));
  orx  g4823(.a(n4863), .b(n4860), .O(n4864));
  orx  g4824(.a(n4864), .b(n4859), .O(n4865));
  andx g4825(.a(pi20), .b(pi19), .O(n4866));
  andx g4826(.a(n4866), .b(pi17), .O(n4867));
  andx g4827(.a(n4867), .b(n3210), .O(n4868));
  andx g4828(.a(n4868), .b(n4136), .O(n4869));
  andx g4829(.a(n3430), .b(n3244), .O(n4870));
  andx g4830(.a(n4870), .b(n3434), .O(n4871));
  orx  g4831(.a(n4871), .b(n4869), .O(n4872));
  andx g4832(.a(n3212), .b(n3180), .O(n4873));
  andx g4833(.a(n4873), .b(n3843), .O(n4874));
  andx g4834(.a(n4874), .b(n3851), .O(n4875));
  andx g4835(.a(n3389), .b(n3195), .O(n4876));
  andx g4836(.a(n3672), .b(n3297), .O(n4877));
  andx g4837(.a(n3199), .b(n1021), .O(n4878));
  andx g4838(.a(n4878), .b(n3203), .O(n4879));
  andx g4839(.a(n4879), .b(n4877), .O(n4880));
  andx g4840(.a(n4880), .b(n4876), .O(n4881));
  orx  g4841(.a(n4881), .b(n4875), .O(n4882));
  orx  g4842(.a(n4882), .b(n4872), .O(n4883));
  orx  g4843(.a(n4883), .b(n4865), .O(n4884));
  orx  g4844(.a(n4884), .b(n4855), .O(n4885));
  andx g4845(.a(n4857), .b(n3781), .O(n4886));
  andx g4846(.a(n3933), .b(n3845), .O(n4887));
  orx  g4847(.a(n4887), .b(n4886), .O(n4888));
  andx g4848(.a(n3214), .b(n92), .O(n4889));
  andx g4849(.a(n4889), .b(n4748), .O(n4890));
  andx g4850(.a(n4890), .b(n3543), .O(n4891));
  andx g4851(.a(n47), .b(n63), .O(n4892));
  andx g4852(.a(n4892), .b(n3624), .O(n4893));
  andx g4853(.a(n3735), .b(n3369), .O(n4894));
  andx g4854(.a(n4894), .b(n4893), .O(n4895));
  andx g4855(.a(n4895), .b(n3385), .O(n4896));
  andx g4856(.a(n4896), .b(n4174), .O(n4897));
  orx  g4857(.a(n4897), .b(n4891), .O(n4898));
  orx  g4858(.a(n4898), .b(n4888), .O(n4899));
  andx g4859(.a(n3664), .b(n3191), .O(n4900));
  andx g4860(.a(n533), .b(n67), .O(n4901));
  andx g4861(.a(n4901), .b(n3297), .O(n4902));
  andx g4862(.a(n3453), .b(n48), .O(n4903));
  andx g4863(.a(n4903), .b(n4902), .O(n4904));
  andx g4864(.a(n4904), .b(n4876), .O(n4905));
  orx  g4865(.a(n4905), .b(n4900), .O(n4906));
  andx g4866(.a(n3788), .b(pi35), .O(n4907));
  andx g4867(.a(n3181), .b(n895), .O(n4908));
  andx g4868(.a(n4908), .b(n3185), .O(n4909));
  andx g4869(.a(n4909), .b(n4907), .O(n4910));
  andx g4870(.a(n3938), .b(n3781), .O(n4911));
  orx  g4871(.a(n4911), .b(n4910), .O(n4912));
  orx  g4872(.a(n4912), .b(n4906), .O(n4913));
  orx  g4873(.a(n4913), .b(n4899), .O(n4914));
  andx g4874(.a(n4867), .b(n3850), .O(n4915));
  andx g4875(.a(n4915), .b(n4768), .O(n4916));
  andx g4876(.a(n3429), .b(n1942), .O(n4917));
  andx g4877(.a(n3253), .b(n303), .O(n4918));
  andx g4878(.a(n4237), .b(n3672), .O(n4919));
  andx g4879(.a(n4919), .b(n4918), .O(n4920));
  andx g4880(.a(n4920), .b(n4917), .O(n4921));
  orx  g4881(.a(n4921), .b(n4916), .O(n4922));
  andx g4882(.a(n3708), .b(n3469), .O(n4923));
  andx g4883(.a(n4923), .b(n45), .O(n4924));
  andx g4884(.a(n4924), .b(n3532), .O(n4925));
  andx g4885(.a(n4925), .b(n4876), .O(n4926));
  andx g4886(.a(n3266), .b(n3186), .O(n4927));
  andx g4887(.a(n4189), .b(n3419), .O(n4928));
  andx g4888(.a(n4928), .b(n4400), .O(n4929));
  andx g4889(.a(n4929), .b(n4927), .O(n4930));
  orx  g4890(.a(n4930), .b(n4926), .O(n4931));
  orx  g4891(.a(n4931), .b(n4922), .O(n4932));
  andx g4892(.a(n3911), .b(n3203), .O(n4933));
  andx g4893(.a(n4933), .b(n3897), .O(n4934));
  andx g4894(.a(n4934), .b(n3478), .O(n4935));
  andx g4895(.a(n3451), .b(n264), .O(n4936));
  andx g4896(.a(n3419), .b(n48), .O(n4937));
  andx g4897(.a(n4937), .b(n4936), .O(n4938));
  andx g4898(.a(n4938), .b(n3789), .O(n4939));
  andx g4899(.a(n4939), .b(n3960), .O(n4940));
  orx  g4900(.a(n4940), .b(n4935), .O(n4941));
  andx g4901(.a(n3871), .b(n3234), .O(n4942));
  andx g4902(.a(n4942), .b(n3708), .O(n4943));
  andx g4903(.a(n4943), .b(n3385), .O(n4944));
  andx g4904(.a(n4944), .b(n3886), .O(n4945));
  andx g4905(.a(n3239), .b(n3221), .O(n4946));
  andx g4906(.a(n3469), .b(n48), .O(n4947));
  andx g4907(.a(n4947), .b(n4946), .O(n4948));
  andx g4908(.a(n4948), .b(n4057), .O(n4949));
  andx g4909(.a(n4949), .b(n3956), .O(n4950));
  orx  g4910(.a(n4950), .b(n4945), .O(n4951));
  orx  g4911(.a(n4951), .b(n4941), .O(n4952));
  orx  g4912(.a(n4952), .b(n4932), .O(n4953));
  orx  g4913(.a(n4953), .b(n4914), .O(n4954));
  orx  g4914(.a(n4954), .b(n4885), .O(n4955));
  andx g4915(.a(n46), .b(n212), .O(n4956));
  andx g4916(.a(n4956), .b(n47), .O(n4957));
  andx g4917(.a(n4957), .b(n45), .O(n4958));
  andx g4918(.a(n4958), .b(n3381), .O(n4959));
  andx g4919(.a(n4748), .b(n3214), .O(n4960));
  andx g4920(.a(n4960), .b(n4959), .O(n4961));
  andx g4921(.a(n3510), .b(n3353), .O(n4962));
  orx  g4922(.a(n4962), .b(n4961), .O(n4963));
  andx g4923(.a(n3449), .b(n43), .O(n4964));
  andx g4924(.a(n3348), .b(n73), .O(n4965));
  andx g4925(.a(n4965), .b(n4134), .O(n4966));
  andx g4926(.a(n4966), .b(n4964), .O(n4967));
  andx g4927(.a(n3374), .b(n2508), .O(n4968));
  andx g4928(.a(n4968), .b(n3441), .O(n4969));
  orx  g4929(.a(n4969), .b(n4967), .O(n4970));
  orx  g4930(.a(n4970), .b(n4963), .O(n4971));
  andx g4931(.a(n3672), .b(n3452), .O(n4972));
  andx g4932(.a(n3253), .b(n3248), .O(n4973));
  andx g4933(.a(n4973), .b(n3203), .O(n4974));
  andx g4934(.a(n4974), .b(n4972), .O(n4975));
  andx g4935(.a(n4975), .b(n3670), .O(n4976));
  andx g4936(.a(n4820), .b(n88), .O(n4977));
  andx g4937(.a(n3290), .b(n67), .O(n4978));
  andx g4938(.a(n3736), .b(n3367), .O(n4979));
  andx g4939(.a(n4979), .b(n4894), .O(n4980));
  andx g4940(.a(n4980), .b(n4978), .O(n4981));
  andx g4941(.a(n4981), .b(n4977), .O(n4982));
  orx  g4942(.a(n4982), .b(n4976), .O(n4983));
  andx g4943(.a(n3320), .b(n3248), .O(n4984));
  andx g4944(.a(n4984), .b(n3267), .O(n4985));
  andx g4945(.a(n4985), .b(n4907), .O(n4986));
  andx g4946(.a(n3824), .b(n3356), .O(n4987));
  orx  g4947(.a(n4987), .b(n4986), .O(n4988));
  orx  g4948(.a(n4988), .b(n4983), .O(n4989));
  orx  g4949(.a(n4989), .b(n4971), .O(n4990));
  andx g4950(.a(n3638), .b(n3475), .O(n4991));
  andx g4951(.a(n48), .b(n303), .O(n4992));
  andx g4952(.a(pi35), .b(n64), .O(n4993));
  andx g4953(.a(n4993), .b(n298), .O(n4994));
  andx g4954(.a(n4994), .b(n4992), .O(n4995));
  andx g4955(.a(n4995), .b(n3431), .O(n4996));
  orx  g4956(.a(n4996), .b(n4991), .O(n4997));
  andx g4957(.a(n1773), .b(n895), .O(n4998));
  andx g4958(.a(n4998), .b(n3708), .O(n4999));
  andx g4959(.a(n4999), .b(n3247), .O(n5000));
  andx g4960(.a(n5000), .b(n3707), .O(n5001));
  andx g4961(.a(n3898), .b(n164), .O(n5002));
  andx g4962(.a(n5002), .b(n4120), .O(n5003));
  andx g4963(.a(n5003), .b(n3374), .O(n5004));
  andx g4964(.a(n5004), .b(n3747), .O(n5005));
  orx  g4965(.a(n5005), .b(n5001), .O(n5006));
  orx  g4966(.a(n5006), .b(n4997), .O(n5007));
  andx g4967(.a(n3422), .b(n73), .O(n5008));
  andx g4968(.a(n5008), .b(n298), .O(n5009));
  andx g4969(.a(n5009), .b(n3421), .O(n5010));
  andx g4970(.a(n5010), .b(n3315), .O(n5011));
  andx g4971(.a(n3420), .b(n65), .O(n5012));
  andx g4972(.a(n5012), .b(n3255), .O(n5013));
  andx g4973(.a(n5013), .b(n3476), .O(n5014));
  andx g4974(.a(n5014), .b(n4964), .O(n5015));
  orx  g4975(.a(n5015), .b(n5011), .O(n5016));
  andx g4976(.a(n3447), .b(n3257), .O(n5017));
  andx g4977(.a(n3232), .b(n3202), .O(n5018));
  andx g4978(.a(n65), .b(n49), .O(n5019));
  andx g4979(.a(n5019), .b(n5018), .O(n5020));
  andx g4980(.a(n5020), .b(n3197), .O(n5021));
  orx  g4981(.a(n5021), .b(n5017), .O(n5022));
  orx  g4982(.a(n5022), .b(n5016), .O(n5023));
  orx  g4983(.a(n5023), .b(n5007), .O(n5024));
  orx  g4984(.a(n5024), .b(n4990), .O(n5025));
  andx g4985(.a(n92), .b(n63), .O(n5026));
  andx g4986(.a(n5026), .b(n3508), .O(n5027));
  andx g4987(.a(n5027), .b(n3560), .O(n5028));
  andx g4988(.a(n1689), .b(n855), .O(n5029));
  andx g4989(.a(n3881), .b(n3672), .O(n5030));
  andx g4990(.a(n5030), .b(n48), .O(n5031));
  andx g4991(.a(n5031), .b(n5029), .O(n5032));
  andx g4992(.a(n5032), .b(n3670), .O(n5033));
  orx  g4993(.a(n5033), .b(n5028), .O(n5034));
  andx g4994(.a(n5027), .b(n3489), .O(n5035));
  andx g4995(.a(n3224), .b(n88), .O(n5036));
  andx g4996(.a(n5036), .b(n3446), .O(n5037));
  orx  g4997(.a(n5037), .b(n5035), .O(n5038));
  orx  g4998(.a(n5038), .b(n5034), .O(n5039));
  andx g4999(.a(n4918), .b(n4154), .O(n5040));
  andx g5000(.a(n5040), .b(n3310), .O(n5041));
  andx g5001(.a(n3199), .b(n2507), .O(n5042));
  andx g5002(.a(n5042), .b(n4822), .O(n5043));
  andx g5003(.a(n5043), .b(n3476), .O(n5044));
  andx g5004(.a(n5044), .b(n4174), .O(n5045));
  orx  g5005(.a(n5045), .b(n5041), .O(n5046));
  andx g5006(.a(n5040), .b(n3583), .O(n5047));
  andx g5007(.a(n4156), .b(n3580), .O(n5048));
  orx  g5008(.a(n5048), .b(n5047), .O(n5049));
  orx  g5009(.a(n5049), .b(n5046), .O(n5050));
  orx  g5010(.a(n5050), .b(n5039), .O(n5051));
  andx g5011(.a(n3898), .b(n1689), .O(n5052));
  andx g5012(.a(n3719), .b(n3367), .O(n5053));
  andx g5013(.a(n5053), .b(n5052), .O(n5054));
  andx g5014(.a(n5054), .b(n4134), .O(n5055));
  andx g5015(.a(n5055), .b(n3366), .O(n5056));
  andx g5016(.a(n3320), .b(n3180), .O(n5057));
  andx g5017(.a(n5057), .b(n3441), .O(n5058));
  orx  g5018(.a(n5058), .b(n5056), .O(n5059));
  andx g5019(.a(n3486), .b(n3471), .O(n5060));
  andx g5020(.a(n3887), .b(n2507), .O(n5061));
  andx g5021(.a(n5061), .b(n3476), .O(n5062));
  andx g5022(.a(n5062), .b(n3392), .O(n5063));
  orx  g5023(.a(n5063), .b(n5060), .O(n5064));
  orx  g5024(.a(n5064), .b(n5059), .O(n5065));
  andx g5025(.a(n4160), .b(n3817), .O(n5066));
  andx g5026(.a(n4861), .b(n3280), .O(n5067));
  orx  g5027(.a(n5067), .b(n5066), .O(n5068));
  andx g5028(.a(n3635), .b(n3478), .O(n5069));
  andx g5029(.a(n5036), .b(n3257), .O(n5070));
  orx  g5030(.a(n5070), .b(n5069), .O(n5071));
  orx  g5031(.a(n5071), .b(n5068), .O(n5072));
  orx  g5032(.a(n5072), .b(n5065), .O(n5073));
  orx  g5033(.a(n5073), .b(n5051), .O(n5074));
  orx  g5034(.a(n5074), .b(n5025), .O(n5075));
  orx  g5035(.a(n5075), .b(n4955), .O(n5076));
  andx g5036(.a(n4851), .b(n4818), .O(n5077));
  andx g5037(.a(pi25), .b(pi26), .O(n5078));
  andx g5038(.a(n5078), .b(n63), .O(n5079));
  andx g5039(.a(n52), .b(pi30), .O(n5080));
  andx g5040(.a(n5080), .b(n4388), .O(n5081));
  andx g5041(.a(n5081), .b(n5079), .O(n5082));
  andx g5042(.a(n5078), .b(n1344), .O(n5083));
  andx g5043(.a(n5083), .b(n4407), .O(n5084));
  orx  g5044(.a(n5084), .b(n5082), .O(n5085));
  andx g5045(.a(n75), .b(pi22), .O(n5086));
  andx g5046(.a(n333), .b(pi29), .O(n5087));
  andx g5047(.a(n5087), .b(n431), .O(n5088));
  andx g5048(.a(n5088), .b(n5086), .O(n5089));
  andx g5049(.a(pi22), .b(n63), .O(n5090));
  andx g5050(.a(n5090), .b(pi30), .O(n5091));
  andx g5051(.a(n5091), .b(n182), .O(n5092));
  orx  g5052(.a(n5092), .b(n5089), .O(n5093));
  orx  g5053(.a(n5093), .b(n5085), .O(n5094));
  orx  g5054(.a(n5094), .b(n5077), .O(n5095));
  andx g5055(.a(n3234), .b(n1688), .O(n5096));
  andx g5056(.a(n5096), .b(n313), .O(n5097));
  andx g5057(.a(n5097), .b(n922), .O(n5098));
  andx g5058(.a(n5098), .b(n3717), .O(n5099));
  andx g5059(.a(n3935), .b(n3842), .O(n5100));
  orx  g5060(.a(n5100), .b(n5099), .O(n5101));
  orx  g5061(.a(n5101), .b(n5095), .O(n5102));
  andx g5062(.a(pi22), .b(pi08), .O(n5103));
  andx g5063(.a(n5103), .b(n230), .O(n5104));
  andx g5064(.a(n199), .b(pi22), .O(n5105));
  andx g5065(.a(n4279), .b(n52), .O(n5106));
  andx g5066(.a(n5106), .b(n5105), .O(n5107));
  orx  g5067(.a(n5107), .b(n5104), .O(n5108));
  andx g5068(.a(pi22), .b(n64), .O(n5109));
  andx g5069(.a(n4388), .b(n437), .O(n5110));
  andx g5070(.a(n5110), .b(n5109), .O(n5111));
  andx g5071(.a(n1344), .b(pi33), .O(n5112));
  andx g5072(.a(n5112), .b(n4407), .O(n5113));
  orx  g5073(.a(n5113), .b(n5111), .O(n5114));
  orx  g5074(.a(n5114), .b(n5108), .O(n5115));
  andx g5075(.a(n431), .b(n110), .O(n5116));
  andx g5076(.a(n5116), .b(n4296), .O(n5117));
  andx g5077(.a(pi22), .b(pi12), .O(n5118));
  andx g5078(.a(n5118), .b(n230), .O(n5119));
  orx  g5079(.a(n5119), .b(n5117), .O(n5120));
  andx g5080(.a(pi22), .b(pi11), .O(n5121));
  andx g5081(.a(n5080), .b(n199), .O(n5122));
  andx g5082(.a(n5122), .b(n5121), .O(n5123));
  andx g5083(.a(n1344), .b(pi32), .O(n5124));
  andx g5084(.a(n5124), .b(n4407), .O(n5125));
  orx  g5085(.a(n5125), .b(n5123), .O(n5126));
  orx  g5086(.a(n5126), .b(n5120), .O(n5127));
  orx  g5087(.a(n5127), .b(n5115), .O(n5128));
  andx g5088(.a(n5080), .b(n4309), .O(n5129));
  andx g5089(.a(n5129), .b(n5079), .O(n5130));
  andx g5090(.a(n5086), .b(n522), .O(n5131));
  orx  g5091(.a(n5131), .b(n5130), .O(n5132));
  andx g5092(.a(pi25), .b(pi09), .O(n5133));
  andx g5093(.a(n5133), .b(n63), .O(n5134));
  andx g5094(.a(pi26), .b(pi08), .O(n5135));
  andx g5095(.a(n5135), .b(n756), .O(n5136));
  andx g5096(.a(n5136), .b(n5134), .O(n5137));
  andx g5097(.a(n5109), .b(n437), .O(n5138));
  andx g5098(.a(n5138), .b(n1815), .O(n5139));
  orx  g5099(.a(n5139), .b(n5137), .O(n5140));
  orx  g5100(.a(n5140), .b(n5132), .O(n5141));
  andx g5101(.a(n5078), .b(pi29), .O(n5142));
  andx g5102(.a(n5142), .b(n3185), .O(n5143));
  andx g5103(.a(n5080), .b(n1815), .O(n5144));
  andx g5104(.a(n5144), .b(n5079), .O(n5145));
  orx  g5105(.a(n5145), .b(n5143), .O(n5146));
  andx g5106(.a(n5122), .b(n1534), .O(n5147));
  andx g5107(.a(n5124), .b(n4629), .O(n5148));
  orx  g5108(.a(n5148), .b(n5147), .O(n5149));
  orx  g5109(.a(n5149), .b(n5146), .O(n5150));
  orx  g5110(.a(n5150), .b(n5141), .O(n5151));
  orx  g5111(.a(n5151), .b(n5128), .O(n5152));
  orx  g5112(.a(n5152), .b(n5102), .O(n5153));
  andx g5113(.a(n43), .b(pi14), .O(n5154));
  andx g5114(.a(n5154), .b(n48), .O(n5155));
  andx g5115(.a(n5155), .b(n3897), .O(n5156));
  andx g5116(.a(n3413), .b(n5156), .O(n5157));
  andx g5117(.a(n3672), .b(n3408), .O(n5158));
  andx g5118(.a(n5158), .b(n4918), .O(n5159));
  andx g5119(.a(n5159), .b(n4917), .O(n5160));
  orx  g5120(.a(n5160), .b(n5157), .O(n5161));
  andx g5121(.a(n3906), .b(n3558), .O(n5162));
  andx g5122(.a(n4960), .b(n3901), .O(n5163));
  orx  g5123(.a(n5163), .b(n5162), .O(n5164));
  orx  g5124(.a(n5164), .b(n5161), .O(n5165));
  andx g5125(.a(n3663), .b(n3183), .O(n5166));
  andx g5126(.a(n3672), .b(n3320), .O(n5167));
  andx g5127(.a(n5167), .b(n3419), .O(n5168));
  andx g5128(.a(n5168), .b(n3742), .O(n5169));
  orx  g5129(.a(n5169), .b(n5166), .O(n5170));
  andx g5130(.a(n301), .b(n48), .O(n5171));
  andx g5131(.a(n5171), .b(n3718), .O(n5172));
  andx g5132(.a(n5172), .b(n3345), .O(n5173));
  andx g5133(.a(n3369), .b(n3202), .O(n5174));
  andx g5134(.a(n3255), .b(n3218), .O(n5175));
  andx g5135(.a(n5175), .b(n5174), .O(n5176));
  andx g5136(.a(n5176), .b(n766), .O(n5177));
  andx g5137(.a(n5177), .b(n3714), .O(n5178));
  orx  g5138(.a(n5178), .b(n5173), .O(n5179));
  orx  g5139(.a(n5179), .b(n5170), .O(n5180));
  orx  g5140(.a(n5180), .b(n5165), .O(n5181));
  orx  g5141(.a(n5181), .b(n5153), .O(n5182));
  andx g5142(.a(n3320), .b(n313), .O(n5183));
  andx g5143(.a(n5183), .b(n3214), .O(n5184));
  andx g5144(.a(n5184), .b(n1439), .O(n5185));
  orx  g5145(.a(n5185), .b(n1521), .O(n5186));
  andx g5146(.a(n4613), .b(n345), .O(n5187));
  andx g5147(.a(n5187), .b(n4686), .O(n5188));
  andx g5148(.a(n5188), .b(n4437), .O(n5189));
  andx g5149(.a(n3577), .b(n644), .O(n5190));
  andx g5150(.a(n5190), .b(n3234), .O(n5191));
  andx g5151(.a(n3367), .b(n675), .O(n5192));
  andx g5152(.a(n3937), .b(n3910), .O(n5193));
  andx g5153(.a(n5193), .b(n5192), .O(n5194));
  andx g5154(.a(n5194), .b(n5191), .O(n5195));
  orx  g5155(.a(n5195), .b(n5189), .O(n5196));
  orx  g5156(.a(n5196), .b(n5186), .O(n5197));
  andx g5157(.a(n3719), .b(n3672), .O(n5198));
  andx g5158(.a(n4608), .b(n3403), .O(n5199));
  andx g5159(.a(n5199), .b(n5198), .O(n5200));
  andx g5160(.a(n5200), .b(n4325), .O(n5201));
  orx  g5161(.a(n5201), .b(n1320), .O(n5202));
  andx g5162(.a(n3734), .b(n5187), .O(n5203));
  andx g5163(.a(n5203), .b(n3404), .O(n5204));
  andx g5164(.a(n4993), .b(n1021), .O(n5205));
  andx g5165(.a(n3194), .b(n1706), .O(n5206));
  andx g5166(.a(n5206), .b(n3231), .O(n5207));
  andx g5167(.a(n5207), .b(n5205), .O(n5208));
  orx  g5168(.a(n5208), .b(n5204), .O(n5209));
  orx  g5169(.a(n5209), .b(n5202), .O(n5210));
  orx  g5170(.a(n5210), .b(n5197), .O(n5211));
  andx g5171(.a(n4608), .b(n3320), .O(n5212));
  andx g5172(.a(n5212), .b(n4288), .O(n5213));
  andx g5173(.a(n5213), .b(n3139), .O(n5214));
  andx g5174(.a(n766), .b(n3270), .O(n5215));
  andx g5175(.a(n5215), .b(n4568), .O(n5216));
  orx  g5176(.a(n5216), .b(n5214), .O(n5217));
  andx g5177(.a(n345), .b(n313), .O(n5218));
  andx g5178(.a(n5218), .b(n4686), .O(n5219));
  andx g5179(.a(n5219), .b(n4685), .O(n5220));
  andx g5180(.a(n3218), .b(n1344), .O(n5221));
  andx g5181(.a(n5221), .b(n3231), .O(n5222));
  andx g5182(.a(n5222), .b(n4728), .O(n5223));
  orx  g5183(.a(n5223), .b(n5220), .O(n5224));
  orx  g5184(.a(n5224), .b(n5217), .O(n5225));
  andx g5185(.a(n4671), .b(n895), .O(n5226));
  andx g5186(.a(n5226), .b(n4471), .O(n5227));
  andx g5187(.a(n3491), .b(n3344), .O(n5228));
  orx  g5188(.a(n5228), .b(n5227), .O(n5229));
  andx g5189(.a(n3416), .b(n73), .O(n5230));
  andx g5190(.a(n4466), .b(n855), .O(n5231));
  andx g5191(.a(n5231), .b(n5230), .O(n5232));
  andx g5192(.a(n3203), .b(n1021), .O(n5233));
  andx g5193(.a(n5233), .b(n3254), .O(n5234));
  andx g5194(.a(n5234), .b(n5232), .O(n5235));
  orx  g5195(.a(n5235), .b(n1264), .O(n5236));
  orx  g5196(.a(n5236), .b(n5229), .O(n5237));
  orx  g5197(.a(n5237), .b(n5225), .O(n5238));
  orx  g5198(.a(n5238), .b(n5211), .O(n5239));
  andx g5199(.a(pi26), .b(pi12), .O(n5240));
  andx g5200(.a(n5240), .b(n756), .O(n5241));
  andx g5201(.a(n5241), .b(n5134), .O(n5242));
  andx g5202(.a(pi12), .b(n63), .O(n5243));
  andx g5203(.a(n5243), .b(n5112), .O(n5244));
  orx  g5204(.a(n5244), .b(n5242), .O(n5245));
  andx g5205(.a(n5078), .b(pi07), .O(n5246));
  andx g5206(.a(n75), .b(pi30), .O(n5247));
  andx g5207(.a(n5247), .b(n4629), .O(n5248));
  andx g5208(.a(n5248), .b(n5246), .O(n5249));
  andx g5209(.a(n4381), .b(n431), .O(n5250));
  andx g5210(.a(n5250), .b(n4296), .O(n5251));
  orx  g5211(.a(n5251), .b(n5249), .O(n5252));
  orx  g5212(.a(n5252), .b(n5245), .O(n5253));
  andx g5213(.a(n5083), .b(n4629), .O(n5254));
  andx g5214(.a(n5243), .b(n5083), .O(n5255));
  orx  g5215(.a(n5255), .b(n5254), .O(n5256));
  andx g5216(.a(n4371), .b(n431), .O(n5257));
  andx g5217(.a(n5257), .b(n4296), .O(n5258));
  andx g5218(.a(n5121), .b(n230), .O(n5259));
  orx  g5219(.a(n5259), .b(n5258), .O(n5260));
  orx  g5220(.a(n5260), .b(n5256), .O(n5261));
  orx  g5221(.a(n5261), .b(n5253), .O(n5262));
  andx g5222(.a(pi25), .b(pi11), .O(n5263));
  andx g5223(.a(pi26), .b(n64), .O(n5264));
  andx g5224(.a(n5264), .b(n5263), .O(n5265));
  andx g5225(.a(n5265), .b(n2713), .O(n5266));
  andx g5226(.a(n5247), .b(n4407), .O(n5267));
  andx g5227(.a(n5267), .b(n5246), .O(n5268));
  orx  g5228(.a(n5268), .b(n5266), .O(n5269));
  andx g5229(.a(n5264), .b(n63), .O(n5270));
  andx g5230(.a(pi07), .b(pi12), .O(n5271));
  andx g5231(.a(n5271), .b(n193), .O(n5272));
  andx g5232(.a(n5272), .b(n5270), .O(n5273));
  andx g5233(.a(n5243), .b(n5124), .O(n5274));
  orx  g5234(.a(n5274), .b(n5273), .O(n5275));
  orx  g5235(.a(n5275), .b(n5269), .O(n5276));
  andx g5236(.a(n5265), .b(n200), .O(n5277));
  andx g5237(.a(n4395), .b(n52), .O(n5278));
  andx g5238(.a(n5278), .b(n5105), .O(n5279));
  orx  g5239(.a(n5279), .b(n5277), .O(n5280));
  andx g5240(.a(n5264), .b(pi07), .O(n5281));
  andx g5241(.a(n4629), .b(n193), .O(n5282));
  andx g5242(.a(n5282), .b(n5281), .O(n5283));
  andx g5243(.a(pi07), .b(pi30), .O(n5284));
  andx g5244(.a(n5284), .b(n229), .O(n5285));
  andx g5245(.a(n5285), .b(n1534), .O(n5286));
  orx  g5246(.a(n5286), .b(n5283), .O(n5287));
  orx  g5247(.a(n5287), .b(n5280), .O(n5288));
  orx  g5248(.a(n5288), .b(n5276), .O(n5289));
  orx  g5249(.a(n5289), .b(n5262), .O(n5290));
  andx g5250(.a(n4608), .b(n3196), .O(n5291));
  andx g5251(.a(n5291), .b(n3941), .O(n5292));
  andx g5252(.a(n5292), .b(n4427), .O(n5293));
  orx  g5253(.a(n5293), .b(n408), .O(n5294));
  andx g5254(.a(n484), .b(n73), .O(n5295));
  andx g5255(.a(n5295), .b(n49), .O(n5296));
  andx g5256(.a(n5296), .b(n4788), .O(n5297));
  andx g5257(.a(n4608), .b(n3856), .O(n5298));
  andx g5258(.a(n5298), .b(n381), .O(n5299));
  andx g5259(.a(n4464), .b(n3241), .O(n5300));
  andx g5260(.a(n5300), .b(n3734), .O(n5301));
  andx g5261(.a(n5301), .b(n5299), .O(n5302));
  orx  g5262(.a(n5302), .b(n5297), .O(n5303));
  orx  g5263(.a(n5303), .b(n5294), .O(n5304));
  andx g5264(.a(n431), .b(pi33), .O(n5305));
  andx g5265(.a(n5305), .b(n4371), .O(n5306));
  andx g5266(.a(n5138), .b(n4309), .O(n5307));
  orx  g5267(.a(n5307), .b(n5306), .O(n5308));
  andx g5268(.a(n5247), .b(n5243), .O(n5309));
  andx g5269(.a(n5309), .b(n5246), .O(n5310));
  andx g5270(.a(n230), .b(n1534), .O(n5311));
  orx  g5271(.a(n5311), .b(n5310), .O(n5312));
  orx  g5272(.a(n5312), .b(n5308), .O(n5313));
  andx g5273(.a(n5296), .b(n4543), .O(n5314));
  andx g5274(.a(n3953), .b(n3708), .O(n5315));
  andx g5275(.a(n2682), .b(n644), .O(n5316));
  andx g5276(.a(n5316), .b(n5315), .O(n5317));
  andx g5277(.a(n45), .b(pi35), .O(n5318));
  andx g5278(.a(n5318), .b(n4431), .O(n5319));
  andx g5279(.a(n5319), .b(n5317), .O(n5320));
  orx  g5280(.a(n5320), .b(n5314), .O(n5321));
  orx  g5281(.a(n5321), .b(n5313), .O(n5322));
  orx  g5282(.a(n5322), .b(n5304), .O(n5323));
  orx  g5283(.a(n5323), .b(n5290), .O(n5324));
  orx  g5284(.a(n5324), .b(n5239), .O(n5325));
  orx  g5285(.a(n5325), .b(n5182), .O(n5326));
  andx g5286(.a(n1831), .b(n299), .O(n5327));
  andx g5287(.a(n5327), .b(n3374), .O(n5328));
  andx g5288(.a(n5328), .b(n3680), .O(n5329));
  andx g5289(.a(n3359), .b(n49), .O(n5330));
  andx g5290(.a(n5330), .b(n3902), .O(n5331));
  orx  g5291(.a(n5331), .b(n5329), .O(n5332));
  andx g5292(.a(n4915), .b(n4251), .O(n5333));
  andx g5293(.a(n3469), .b(n3261), .O(n5334));
  andx g5294(.a(n5334), .b(n45), .O(n5335));
  andx g5295(.a(n5335), .b(n3588), .O(n5336));
  andx g5296(.a(n5336), .b(n3499), .O(n5337));
  orx  g5297(.a(n5337), .b(n5333), .O(n5338));
  orx  g5298(.a(n5338), .b(n5332), .O(n5339));
  andx g5299(.a(n3272), .b(n3218), .O(n5340));
  andx g5300(.a(n5340), .b(n3480), .O(n5341));
  andx g5301(.a(n5341), .b(n4927), .O(n5342));
  andx g5302(.a(n3246), .b(n3232), .O(n5343));
  andx g5303(.a(n4892), .b(n3261), .O(n5344));
  andx g5304(.a(n5344), .b(n45), .O(n5345));
  andx g5305(.a(n5345), .b(n5343), .O(n5346));
  andx g5306(.a(n5346), .b(n3295), .O(n5347));
  orx  g5307(.a(n5347), .b(n5342), .O(n5348));
  andx g5308(.a(n3246), .b(n87), .O(n5349));
  andx g5309(.a(n3856), .b(n3203), .O(n5350));
  andx g5310(.a(n5350), .b(n313), .O(n5351));
  andx g5311(.a(n5351), .b(n5349), .O(n5352));
  andx g5312(.a(n5352), .b(n4876), .O(n5353));
  andx g5313(.a(n4851), .b(n3893), .O(n5354));
  orx  g5314(.a(n5354), .b(n5353), .O(n5355));
  orx  g5315(.a(n5355), .b(n5348), .O(n5356));
  orx  g5316(.a(n5356), .b(n5339), .O(n5357));
  andx g5317(.a(n3902), .b(n4959), .O(n5358));
  andx g5318(.a(n4939), .b(n3956), .O(n5359));
  orx  g5319(.a(n5359), .b(n5358), .O(n5360));
  andx g5320(.a(n4161), .b(n4868), .O(n5361));
  andx g5321(.a(n4995), .b(n4870), .O(n5362));
  orx  g5322(.a(n5362), .b(n5361), .O(n5363));
  orx  g5323(.a(n5363), .b(n5360), .O(n5364));
  andx g5324(.a(n895), .b(n63), .O(n5365));
  andx g5325(.a(n3735), .b(n2832), .O(n5366));
  andx g5326(.a(n5366), .b(n3734), .O(n5367));
  andx g5327(.a(n5367), .b(n5365), .O(n5368));
  andx g5328(.a(n5368), .b(n4821), .O(n5369));
  andx g5329(.a(n4088), .b(n3406), .O(n5370));
  andx g5330(.a(n5370), .b(n4822), .O(n5371));
  andx g5331(.a(n5371), .b(n3687), .O(n5372));
  andx g5332(.a(n5372), .b(n4977), .O(n5373));
  orx  g5333(.a(n5373), .b(n5369), .O(n5374));
  andx g5334(.a(n4934), .b(n3638), .O(n5375));
  andx g5335(.a(n4949), .b(n3960), .O(n5376));
  orx  g5336(.a(n5376), .b(n5375), .O(n5377));
  orx  g5337(.a(n5377), .b(n5374), .O(n5378));
  orx  g5338(.a(n5378), .b(n5364), .O(n5379));
  orx  g5339(.a(n5379), .b(n5357), .O(n5380));
  andx g5340(.a(n3382), .b(n65), .O(n5381));
  andx g5341(.a(n5381), .b(n4497), .O(n5382));
  andx g5342(.a(n5382), .b(n3385), .O(n5383));
  andx g5343(.a(n5383), .b(n3295), .O(n5384));
  andx g5344(.a(n4607), .b(n3736), .O(n5385));
  andx g5345(.a(n5385), .b(n3290), .O(n5386));
  andx g5346(.a(n5386), .b(n1209), .O(n5387));
  andx g5347(.a(n5387), .b(n3539), .O(n5388));
  orx  g5348(.a(n5388), .b(n5384), .O(n5389));
  andx g5349(.a(n5040), .b(n3703), .O(n5390));
  andx g5350(.a(n3708), .b(n3406), .O(n5391));
  andx g5351(.a(n5391), .b(n2507), .O(n5392));
  andx g5352(.a(n5392), .b(n3687), .O(n5393));
  andx g5353(.a(n5393), .b(n3742), .O(n5394));
  orx  g5354(.a(n5394), .b(n5390), .O(n5395));
  orx  g5355(.a(n5395), .b(n5389), .O(n5396));
  andx g5356(.a(n3654), .b(n3510), .O(n5397));
  andx g5357(.a(n3406), .b(n644), .O(n5398));
  andx g5358(.a(n5398), .b(n3203), .O(n5399));
  andx g5359(.a(n5399), .b(n3386), .O(n5400));
  andx g5360(.a(n5400), .b(n3717), .O(n5401));
  orx  g5361(.a(n5401), .b(n5397), .O(n5402));
  andx g5362(.a(n5330), .b(n4960), .O(n5403));
  andx g5363(.a(n4924), .b(n3671), .O(n5404));
  andx g5364(.a(n5404), .b(n3670), .O(n5405));
  orx  g5365(.a(n5405), .b(n5403), .O(n5406));
  orx  g5366(.a(n5406), .b(n5402), .O(n5407));
  orx  g5367(.a(n5407), .b(n5396), .O(n5408));
  andx g5368(.a(n4236), .b(n3882), .O(n5409));
  andx g5369(.a(n5409), .b(n3880), .O(n5410));
  andx g5370(.a(n5410), .b(n3879), .O(n5411));
  andx g5371(.a(n3715), .b(n3257), .O(n5412));
  orx  g5372(.a(n5412), .b(n5411), .O(n5413));
  andx g5373(.a(n3913), .b(n3822), .O(n5414));
  andx g5374(.a(n3446), .b(n3263), .O(n5415));
  orx  g5375(.a(n5415), .b(n5414), .O(n5416));
  orx  g5376(.a(n5416), .b(n5413), .O(n5417));
  andx g5377(.a(n5040), .b(n3798), .O(n5418));
  andx g5378(.a(n3736), .b(n3255), .O(n5419));
  andx g5379(.a(n5419), .b(n4894), .O(n5420));
  andx g5380(.a(n5420), .b(n3476), .O(n5421));
  andx g5381(.a(n5421), .b(n3733), .O(n5422));
  orx  g5382(.a(n5422), .b(n5418), .O(n5423));
  andx g5383(.a(n3406), .b(n153), .O(n5424));
  andx g5384(.a(n5424), .b(n3203), .O(n5425));
  andx g5385(.a(n5425), .b(n3271), .O(n5426));
  andx g5386(.a(n5426), .b(n3198), .O(n5427));
  andx g5387(.a(n5156), .b(n3387), .O(n5428));
  orx  g5388(.a(n5428), .b(n5427), .O(n5429));
  orx  g5389(.a(n5429), .b(n5423), .O(n5430));
  orx  g5390(.a(n5430), .b(n5417), .O(n5431));
  orx  g5391(.a(n5431), .b(n5408), .O(n5432));
  orx  g5392(.a(n5432), .b(n5380), .O(n5433));
  orx  g5393(.a(n5433), .b(n5326), .O(n5434));
  orx  g5394(.a(n5434), .b(n5076), .O(n5435));
  orx  g5395(.a(n5435), .b(n4817), .O(n5436));
  orx  g5396(.a(n5436), .b(n4277), .O(n5437));
  orx  g5397(.a(n5437), .b(n4086), .O(po2));
endmodule


