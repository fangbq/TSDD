// Benchmark "sqrt32" written by ABC on Fri Feb  7 13:47:56 2014

module sqrt32 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
    n76, n77, n78, n80, n81, n83, n84, n85, n87, n88, n89, n91, n92, n93,
    n94, n95, n96, n98, n99, n101, n102, n104, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n121, n122,
    n124, n125, n127, n128, n129, n131, n133, n134, n135, n136, n137, n138,
    n140, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295;
  bufx g0000(.A(n918), .O(n48));
  bufx g0001(.A(n918), .O(n49));
  bufx g0002(.A(n403), .O(n50));
  bufx g0003(.A(n403), .O(n51));
  bufx g0004(.A(n527), .O(n52));
  bufx g0005(.A(n527), .O(n53));
  bufx g0006(.A(n831), .O(n54));
  bufx g0007(.A(n831), .O(n55));
  bufx g0008(.A(n742), .O(n56));
  bufx g0009(.A(n742), .O(n57));
  bufx g0010(.A(n742), .O(n58));
  bufx g0011(.A(n1259), .O(n59));
  bufx g0012(.A(n1259), .O(n60));
  bufx g0013(.A(n1259), .O(n61));
  bufx g0014(.A(n1063), .O(n62));
  bufx g0015(.A(n1063), .O(n63));
  bufx g0016(.A(n1063), .O(n64));
  bufx g0017(.A(n84), .O(n65));
  bufx g0018(.A(n84), .O(n66));
  bufx g0019(.A(n84), .O(n67));
  bufx g0020(.A(n84), .O(n68));
  bufx g0021(.A(n1218), .O(n69));
  bufx g0022(.A(n1218), .O(n70));
  bufx g0023(.A(n1218), .O(n71));
  bufx g0024(.A(n636), .O(n72));
  bufx g0025(.A(n636), .O(n73));
  bufx g0026(.A(n96), .O(n74));
  bufx g0027(.A(n96), .O(n75));
  bufx g0028(.A(n96), .O(n76));
  bufx g0029(.A(n96), .O(n77));
  bufx g0030(.A(n843), .O(n78));
  bufx g0031(.A(n843), .O(po06));
  bufx g0032(.A(n843), .O(n80));
  bufx g0033(.A(n415), .O(n81));
  bufx g0034(.A(n415), .O(po02));
  bufx g0035(.A(n415), .O(n83));
  invx g0036(.A(n1129), .O(n84));
  invx g0037(.A(n84), .O(n85));
  invx g0038(.A(n84), .O(po10));
  invx g0039(.A(n84), .O(n87));
  invx g0040(.A(n1219), .O(n88));
  invx g0041(.A(n88), .O(n89));
  invx g0042(.A(n88), .O(po12));
  invx g0043(.A(n88), .O(n91));
  bufx g0044(.A(n282), .O(n92));
  bufx g0045(.A(n282), .O(n93));
  bufx g0046(.A(n1266), .O(n94));
  bufx g0047(.A(n1266), .O(n95));
  invx g0048(.A(n1006), .O(n96));
  invx g0049(.A(n96), .O(po08));
  invx g0050(.A(n96), .O(n98));
  bufx g0051(.A(n751), .O(n99));
  bufx g0052(.A(n751), .O(po05));
  bufx g0053(.A(n751), .O(n101));
  bufx g0054(.A(n536), .O(n102));
  bufx g0055(.A(n536), .O(po03));
  bufx g0056(.A(n536), .O(n104));
  bufx g0057(.A(n1250), .O(po13));
  bufx g0058(.A(n1250), .O(n106));
  bufx g0059(.A(n1250), .O(n107));
  bufx g0060(.A(po11), .O(n108));
  bufx g0061(.A(po11), .O(n109));
  bufx g0062(.A(po11), .O(n110));
  invx g0063(.A(n1168), .O(n111));
  invx g0064(.A(n111), .O(n112));
  invx g0065(.A(n111), .O(n113));
  invx g0066(.A(n111), .O(n114));
  invx g0067(.A(n1241), .O(n115));
  invx g0068(.A(n115), .O(n116));
  invx g0069(.A(n115), .O(n117));
  invx g0070(.A(n115), .O(n118));
  bufx g0071(.A(n283), .O(n119));
  bufx g0072(.A(n283), .O(po01));
  bufx g0073(.A(n283), .O(n121));
  bufx g0074(.A(n648), .O(n122));
  bufx g0075(.A(n648), .O(po04));
  bufx g0076(.A(n648), .O(n124));
  bufx g0077(.A(n1072), .O(n125));
  bufx g0078(.A(n1072), .O(po09));
  bufx g0079(.A(n1072), .O(n127));
  bufx g0080(.A(n927), .O(n128));
  bufx g0081(.A(n927), .O(n129));
  bufx g0082(.A(n927), .O(po07));
  invx g0083(.A(n1268), .O(n131));
  invx g0084(.A(n131), .O(po15));
  invx g0085(.A(n131), .O(n133));
  invx g0086(.A(n131), .O(n134));
  invx g0087(.A(n131), .O(n135));
  invx g0088(.A(n1276), .O(n136));
  invx g0089(.A(n136), .O(n137));
  invx g0090(.A(n136), .O(n138));
  invx g0091(.A(n136), .O(po14));
  invx g0092(.A(n136), .O(n140));
  orx  g0093(.A(n146), .B(n142), .O(po00));
  orx  g0094(.A(n145), .B(n143), .O(n142));
  invx g0095(.A(n144), .O(n143));
  orx  g0096(.A(n287), .B(n92), .O(n144));
  andx g0097(.A(n153), .B(n278), .O(n145));
  orx  g0098(.A(n149), .B(n147), .O(n146));
  andx g0099(.A(n148), .B(n134), .O(n147));
  andx g0100(.A(n296), .B(n288), .O(n148));
  andx g0101(.A(n150), .B(n61), .O(n149));
  orx  g0102(.A(n278), .B(n151), .O(n150));
  orx  g0103(.A(n153), .B(n152), .O(n151));
  andx g0104(.A(n295), .B(n288), .O(n152));
  invx g0105(.A(n154), .O(n153));
  orx  g0106(.A(n156), .B(n155), .O(n154));
  andx g0107(.A(n273), .B(n158), .O(n155));
  andx g0108(.A(n157), .B(po14), .O(n156));
  orx  g0109(.A(n273), .B(n158), .O(n157));
  orx  g0110(.A(n160), .B(n159), .O(n158));
  andx g0111(.A(n268), .B(n162), .O(n159));
  andx g0112(.A(n161), .B(po13), .O(n160));
  orx  g0113(.A(n268), .B(n162), .O(n161));
  orx  g0114(.A(n164), .B(n163), .O(n162));
  andx g0115(.A(n263), .B(n166), .O(n163));
  andx g0116(.A(n165), .B(n89), .O(n164));
  orx  g0117(.A(n263), .B(n166), .O(n165));
  orx  g0118(.A(n168), .B(n167), .O(n166));
  andx g0119(.A(n258), .B(n170), .O(n167));
  andx g0120(.A(n169), .B(po11), .O(n168));
  orx  g0121(.A(n258), .B(n170), .O(n169));
  orx  g0122(.A(n172), .B(n171), .O(n170));
  andx g0123(.A(n253), .B(n174), .O(n171));
  andx g0124(.A(n173), .B(n85), .O(n172));
  orx  g0125(.A(n253), .B(n174), .O(n173));
  orx  g0126(.A(n176), .B(n175), .O(n174));
  andx g0127(.A(n248), .B(n178), .O(n175));
  andx g0128(.A(n177), .B(n125), .O(n176));
  orx  g0129(.A(n248), .B(n178), .O(n177));
  orx  g0130(.A(n180), .B(n179), .O(n178));
  andx g0131(.A(n243), .B(n182), .O(n179));
  andx g0132(.A(n181), .B(n1006), .O(n180));
  orx  g0133(.A(n243), .B(n182), .O(n181));
  orx  g0134(.A(n184), .B(n183), .O(n182));
  andx g0135(.A(n238), .B(n186), .O(n183));
  andx g0136(.A(n185), .B(n927), .O(n184));
  orx  g0137(.A(n238), .B(n186), .O(n185));
  orx  g0138(.A(n188), .B(n187), .O(n186));
  andx g0139(.A(n233), .B(n190), .O(n187));
  andx g0140(.A(n189), .B(n80), .O(n188));
  orx  g0141(.A(n233), .B(n190), .O(n189));
  orx  g0142(.A(n192), .B(n191), .O(n190));
  andx g0143(.A(n228), .B(n194), .O(n191));
  andx g0144(.A(n193), .B(n751), .O(n192));
  orx  g0145(.A(n228), .B(n194), .O(n193));
  orx  g0146(.A(n196), .B(n195), .O(n194));
  andx g0147(.A(n223), .B(n198), .O(n195));
  andx g0148(.A(n197), .B(n648), .O(n196));
  orx  g0149(.A(n223), .B(n198), .O(n197));
  orx  g0150(.A(n200), .B(n199), .O(n198));
  andx g0151(.A(n218), .B(n202), .O(n199));
  andx g0152(.A(n201), .B(n536), .O(n200));
  orx  g0153(.A(n218), .B(n202), .O(n201));
  orx  g0154(.A(n204), .B(n203), .O(n202));
  andx g0155(.A(n213), .B(n206), .O(n203));
  andx g0156(.A(n205), .B(n415), .O(n204));
  orx  g0157(.A(n213), .B(n206), .O(n205));
  orx  g0158(.A(n208), .B(n207), .O(n206));
  andx g0159(.A(n212), .B(n119), .O(n207));
  andx g0160(.A(n211), .B(n209), .O(n208));
  invx g0161(.A(n210), .O(n209));
  orx  g0162(.A(pi01), .B(pi00), .O(n210));
  orx  g0163(.A(n212), .B(po01), .O(n211));
  xorx g0164(.A(n92), .B(pi02), .O(n212));
  invx g0165(.A(n214), .O(n213));
  orx  g0166(.A(n216), .B(n215), .O(n214));
  andx g0167(.A(n412), .B(n119), .O(n215));
  andx g0168(.A(pi03), .B(n217), .O(n216));
  orx  g0169(.A(n93), .B(pi02), .O(n217));
  invx g0170(.A(n219), .O(n218));
  orx  g0171(.A(n221), .B(n220), .O(n219));
  andx g0172(.A(n407), .B(n119), .O(n220));
  andx g0173(.A(n410), .B(n222), .O(n221));
  orx  g0174(.A(n282), .B(n409), .O(n222));
  invx g0175(.A(n224), .O(n223));
  orx  g0176(.A(n226), .B(n225), .O(n224));
  andx g0177(.A(n397), .B(po01), .O(n225));
  andx g0178(.A(n227), .B(n399), .O(n226));
  orx  g0179(.A(n92), .B(n404), .O(n227));
  invx g0180(.A(n229), .O(n228));
  orx  g0181(.A(n231), .B(n230), .O(n229));
  andx g0182(.A(n388), .B(n121), .O(n230));
  andx g0183(.A(n232), .B(n390), .O(n231));
  orx  g0184(.A(n93), .B(n394), .O(n232));
  invx g0185(.A(n234), .O(n233));
  orx  g0186(.A(n236), .B(n235), .O(n234));
  andx g0187(.A(n379), .B(n283), .O(n235));
  andx g0188(.A(n237), .B(n381), .O(n236));
  orx  g0189(.A(n93), .B(n385), .O(n237));
  invx g0190(.A(n239), .O(n238));
  orx  g0191(.A(n241), .B(n240), .O(n239));
  andx g0192(.A(n370), .B(po01), .O(n240));
  andx g0193(.A(n242), .B(n372), .O(n241));
  orx  g0194(.A(n92), .B(n376), .O(n242));
  invx g0195(.A(n244), .O(n243));
  orx  g0196(.A(n246), .B(n245), .O(n244));
  andx g0197(.A(n361), .B(n121), .O(n245));
  andx g0198(.A(n247), .B(n363), .O(n246));
  orx  g0199(.A(n93), .B(n367), .O(n247));
  invx g0200(.A(n249), .O(n248));
  orx  g0201(.A(n251), .B(n250), .O(n249));
  andx g0202(.A(n352), .B(n121), .O(n250));
  andx g0203(.A(n252), .B(n354), .O(n251));
  orx  g0204(.A(n282), .B(n358), .O(n252));
  invx g0205(.A(n254), .O(n253));
  orx  g0206(.A(n256), .B(n255), .O(n254));
  andx g0207(.A(n343), .B(po01), .O(n255));
  andx g0208(.A(n257), .B(n345), .O(n256));
  orx  g0209(.A(n92), .B(n349), .O(n257));
  invx g0210(.A(n259), .O(n258));
  orx  g0211(.A(n261), .B(n260), .O(n259));
  andx g0212(.A(n334), .B(n121), .O(n260));
  andx g0213(.A(n262), .B(n336), .O(n261));
  orx  g0214(.A(n93), .B(n340), .O(n262));
  invx g0215(.A(n264), .O(n263));
  orx  g0216(.A(n266), .B(n265), .O(n264));
  andx g0217(.A(n325), .B(n119), .O(n265));
  andx g0218(.A(n267), .B(n327), .O(n266));
  orx  g0219(.A(n282), .B(n331), .O(n267));
  invx g0220(.A(n269), .O(n268));
  orx  g0221(.A(n271), .B(n270), .O(n269));
  andx g0222(.A(n316), .B(po01), .O(n270));
  andx g0223(.A(n272), .B(n318), .O(n271));
  orx  g0224(.A(n92), .B(n322), .O(n272));
  invx g0225(.A(n274), .O(n273));
  orx  g0226(.A(n276), .B(n275), .O(n274));
  andx g0227(.A(n307), .B(n121), .O(n275));
  andx g0228(.A(n277), .B(n309), .O(n276));
  orx  g0229(.A(n93), .B(n313), .O(n277));
  orx  g0230(.A(n280), .B(n279), .O(n278));
  andx g0231(.A(n297), .B(po01), .O(n279));
  andx g0232(.A(n281), .B(n299), .O(n280));
  orx  g0233(.A(n282), .B(n304), .O(n281));
  invx g0234(.A(n119), .O(n282));
  orx  g0235(.A(n414), .B(n284), .O(n283));
  orx  g0236(.A(n286), .B(n285), .O(n284));
  andx g0237(.A(n429), .B(n424), .O(n285));
  andx g0238(.A(n294), .B(n287), .O(n286));
  orx  g0239(.A(n293), .B(n288), .O(n287));
  orx  g0240(.A(n291), .B(n289), .O(n288));
  invx g0241(.A(n290), .O(n289));
  orx  g0242(.A(n431), .B(n51), .O(n290));
  andx g0243(.A(n292), .B(n432), .O(n291));
  orx  g0244(.A(n50), .B(n437), .O(n292));
  xorx g0245(.A(n296), .B(n61), .O(n293));
  orx  g0246(.A(n295), .B(n60), .O(n294));
  invx g0247(.A(n296), .O(n295));
  orx  g0248(.A(n305), .B(n297), .O(n296));
  invx g0249(.A(n298), .O(n297));
  orx  g0250(.A(n304), .B(n299), .O(n298));
  orx  g0251(.A(n302), .B(n300), .O(n299));
  invx g0252(.A(n301), .O(n300));
  orx  g0253(.A(n440), .B(n50), .O(n301));
  andx g0254(.A(n303), .B(n441), .O(n302));
  orx  g0255(.A(n51), .B(n445), .O(n303));
  xorx g0256(.A(n306), .B(n95), .O(n304));
  andx g0257(.A(n306), .B(n140), .O(n305));
  orx  g0258(.A(n314), .B(n307), .O(n306));
  invx g0259(.A(n308), .O(n307));
  orx  g0260(.A(n313), .B(n309), .O(n308));
  orx  g0261(.A(n311), .B(n310), .O(n309));
  andx g0262(.A(n449), .B(n81), .O(n310));
  andx g0263(.A(n312), .B(n451), .O(n311));
  orx  g0264(.A(n51), .B(n455), .O(n312));
  xorx g0265(.A(n315), .B(n118), .O(n313));
  andx g0266(.A(n315), .B(n106), .O(n314));
  orx  g0267(.A(n323), .B(n316), .O(n315));
  invx g0268(.A(n317), .O(n316));
  orx  g0269(.A(n322), .B(n318), .O(n317));
  orx  g0270(.A(n320), .B(n319), .O(n318));
  andx g0271(.A(n458), .B(po02), .O(n319));
  andx g0272(.A(n321), .B(n460), .O(n320));
  orx  g0273(.A(n50), .B(n464), .O(n321));
  xorx g0274(.A(n324), .B(n69), .O(n322));
  andx g0275(.A(n324), .B(n89), .O(n323));
  orx  g0276(.A(n332), .B(n325), .O(n324));
  invx g0277(.A(n326), .O(n325));
  orx  g0278(.A(n331), .B(n327), .O(n326));
  orx  g0279(.A(n329), .B(n328), .O(n327));
  andx g0280(.A(n467), .B(n83), .O(n328));
  andx g0281(.A(n330), .B(n469), .O(n329));
  orx  g0282(.A(n51), .B(n473), .O(n330));
  xorx g0283(.A(n333), .B(n112), .O(n331));
  andx g0284(.A(n333), .B(n108), .O(n332));
  orx  g0285(.A(n341), .B(n334), .O(n333));
  invx g0286(.A(n335), .O(n334));
  orx  g0287(.A(n340), .B(n336), .O(n335));
  orx  g0288(.A(n338), .B(n337), .O(n336));
  andx g0289(.A(n476), .B(n83), .O(n337));
  andx g0290(.A(n339), .B(n478), .O(n338));
  orx  g0291(.A(n403), .B(n482), .O(n339));
  xorx g0292(.A(n342), .B(n68), .O(n340));
  andx g0293(.A(n342), .B(n85), .O(n341));
  orx  g0294(.A(n350), .B(n343), .O(n342));
  invx g0295(.A(n344), .O(n343));
  orx  g0296(.A(n349), .B(n345), .O(n344));
  orx  g0297(.A(n347), .B(n346), .O(n345));
  andx g0298(.A(n485), .B(n81), .O(n346));
  andx g0299(.A(n348), .B(n487), .O(n347));
  orx  g0300(.A(n50), .B(n491), .O(n348));
  xorx g0301(.A(n351), .B(n64), .O(n349));
  andx g0302(.A(n351), .B(n125), .O(n350));
  orx  g0303(.A(n359), .B(n352), .O(n351));
  invx g0304(.A(n353), .O(n352));
  orx  g0305(.A(n358), .B(n354), .O(n353));
  orx  g0306(.A(n356), .B(n355), .O(n354));
  andx g0307(.A(n494), .B(po02), .O(n355));
  andx g0308(.A(n357), .B(n496), .O(n356));
  orx  g0309(.A(n51), .B(n500), .O(n357));
  xorx g0310(.A(n360), .B(n75), .O(n358));
  andx g0311(.A(n360), .B(n98), .O(n359));
  orx  g0312(.A(n368), .B(n361), .O(n360));
  invx g0313(.A(n362), .O(n361));
  orx  g0314(.A(n367), .B(n363), .O(n362));
  orx  g0315(.A(n365), .B(n364), .O(n363));
  andx g0316(.A(n503), .B(n83), .O(n364));
  andx g0317(.A(n366), .B(n505), .O(n365));
  orx  g0318(.A(n403), .B(n509), .O(n366));
  xorx g0319(.A(n369), .B(n48), .O(n367));
  andx g0320(.A(n369), .B(n128), .O(n368));
  orx  g0321(.A(n377), .B(n370), .O(n369));
  invx g0322(.A(n371), .O(n370));
  orx  g0323(.A(n376), .B(n372), .O(n371));
  orx  g0324(.A(n374), .B(n373), .O(n372));
  andx g0325(.A(n512), .B(po02), .O(n373));
  andx g0326(.A(n375), .B(n514), .O(n374));
  orx  g0327(.A(n50), .B(n518), .O(n375));
  xorx g0328(.A(n378), .B(n831), .O(n376));
  andx g0329(.A(n378), .B(n843), .O(n377));
  orx  g0330(.A(n386), .B(n379), .O(n378));
  invx g0331(.A(n380), .O(n379));
  orx  g0332(.A(n385), .B(n381), .O(n380));
  orx  g0333(.A(n383), .B(n382), .O(n381));
  andx g0334(.A(n521), .B(n81), .O(n382));
  andx g0335(.A(n384), .B(n523), .O(n383));
  orx  g0336(.A(n51), .B(n528), .O(n384));
  xorx g0337(.A(n387), .B(n58), .O(n385));
  andx g0338(.A(n387), .B(n99), .O(n386));
  orx  g0339(.A(n395), .B(n388), .O(n387));
  invx g0340(.A(n389), .O(n388));
  orx  g0341(.A(n394), .B(n390), .O(n389));
  orx  g0342(.A(n392), .B(n391), .O(n390));
  andx g0343(.A(n531), .B(po02), .O(n391));
  andx g0344(.A(n534), .B(n393), .O(n392));
  orx  g0345(.A(n403), .B(n533), .O(n393));
  xorx g0346(.A(n396), .B(n73), .O(n394));
  andx g0347(.A(n396), .B(n122), .O(n395));
  orx  g0348(.A(n405), .B(n397), .O(n396));
  invx g0349(.A(n398), .O(n397));
  orx  g0350(.A(n404), .B(n399), .O(n398));
  orx  g0351(.A(n401), .B(n400), .O(n399));
  andx g0352(.A(n1294), .B(n83), .O(n400));
  andx g0353(.A(pi05), .B(n402), .O(n401));
  orx  g0354(.A(n50), .B(pi04), .O(n402));
  invx g0355(.A(n83), .O(n403));
  xorx g0356(.A(n406), .B(n52), .O(n404));
  andx g0357(.A(n406), .B(n102), .O(n405));
  orx  g0358(.A(n411), .B(n407), .O(n406));
  invx g0359(.A(n408), .O(n407));
  orx  g0360(.A(n410), .B(n409), .O(n408));
  xorx g0361(.A(n81), .B(n413), .O(n409));
  xorx g0362(.A(po02), .B(pi04), .O(n410));
  andx g0363(.A(n412), .B(n83), .O(n411));
  invx g0364(.A(n413), .O(n412));
  orx  g0365(.A(pi03), .B(pi02), .O(n413));
  andx g0366(.A(n422), .B(n81), .O(n414));
  orx  g0367(.A(n420), .B(n416), .O(n415));
  orx  g0368(.A(n418), .B(n417), .O(n416));
  andx g0369(.A(n546), .B(n541), .O(n417));
  andx g0370(.A(n419), .B(n423), .O(n418));
  orx  g0371(.A(n430), .B(n61), .O(n419));
  andx g0372(.A(n421), .B(po03), .O(n420));
  invx g0373(.A(n540), .O(n421));
  invx g0374(.A(n423), .O(n422));
  orx  g0375(.A(n429), .B(n424), .O(n423));
  orx  g0376(.A(n427), .B(n425), .O(n424));
  invx g0377(.A(n426), .O(n425));
  orx  g0378(.A(n549), .B(n53), .O(n426));
  andx g0379(.A(n428), .B(n550), .O(n427));
  orx  g0380(.A(n52), .B(n555), .O(n428));
  xorx g0381(.A(n430), .B(po15), .O(n429));
  andx g0382(.A(n438), .B(n431), .O(n430));
  orx  g0383(.A(n437), .B(n432), .O(n431));
  orx  g0384(.A(n435), .B(n433), .O(n432));
  invx g0385(.A(n434), .O(n433));
  orx  g0386(.A(n558), .B(n527), .O(n434));
  andx g0387(.A(n436), .B(n559), .O(n435));
  orx  g0388(.A(n53), .B(n563), .O(n436));
  xorx g0389(.A(n439), .B(n137), .O(n437));
  orx  g0390(.A(n439), .B(n95), .O(n438));
  andx g0391(.A(n446), .B(n440), .O(n439));
  orx  g0392(.A(n445), .B(n441), .O(n440));
  orx  g0393(.A(n443), .B(n442), .O(n441));
  andx g0394(.A(n567), .B(n104), .O(n442));
  andx g0395(.A(n444), .B(n569), .O(n443));
  orx  g0396(.A(n53), .B(n573), .O(n444));
  xorx g0397(.A(n448), .B(n117), .O(n445));
  invx g0398(.A(n447), .O(n446));
  andx g0399(.A(n448), .B(n107), .O(n447));
  orx  g0400(.A(n456), .B(n449), .O(n448));
  invx g0401(.A(n450), .O(n449));
  orx  g0402(.A(n455), .B(n451), .O(n450));
  orx  g0403(.A(n453), .B(n452), .O(n451));
  andx g0404(.A(n576), .B(n104), .O(n452));
  andx g0405(.A(n454), .B(n578), .O(n453));
  orx  g0406(.A(n52), .B(n582), .O(n454));
  xorx g0407(.A(n457), .B(n88), .O(n455));
  andx g0408(.A(n457), .B(n89), .O(n456));
  orx  g0409(.A(n465), .B(n458), .O(n457));
  invx g0410(.A(n459), .O(n458));
  orx  g0411(.A(n464), .B(n460), .O(n459));
  orx  g0412(.A(n462), .B(n461), .O(n460));
  andx g0413(.A(n585), .B(n102), .O(n461));
  andx g0414(.A(n463), .B(n587), .O(n462));
  orx  g0415(.A(n53), .B(n591), .O(n463));
  xorx g0416(.A(n466), .B(n114), .O(n464));
  andx g0417(.A(n466), .B(n109), .O(n465));
  orx  g0418(.A(n474), .B(n467), .O(n466));
  invx g0419(.A(n468), .O(n467));
  orx  g0420(.A(n473), .B(n469), .O(n468));
  orx  g0421(.A(n471), .B(n470), .O(n469));
  andx g0422(.A(n594), .B(po03), .O(n470));
  andx g0423(.A(n472), .B(n596), .O(n471));
  orx  g0424(.A(n527), .B(n600), .O(n472));
  xorx g0425(.A(n475), .B(n67), .O(n473));
  andx g0426(.A(n475), .B(n87), .O(n474));
  orx  g0427(.A(n483), .B(n476), .O(n475));
  invx g0428(.A(n477), .O(n476));
  orx  g0429(.A(n482), .B(n478), .O(n477));
  orx  g0430(.A(n480), .B(n479), .O(n478));
  andx g0431(.A(n603), .B(n104), .O(n479));
  andx g0432(.A(n481), .B(n605), .O(n480));
  orx  g0433(.A(n52), .B(n609), .O(n481));
  xorx g0434(.A(n484), .B(n63), .O(n482));
  andx g0435(.A(n484), .B(n127), .O(n483));
  orx  g0436(.A(n492), .B(n485), .O(n484));
  invx g0437(.A(n486), .O(n485));
  orx  g0438(.A(n491), .B(n487), .O(n486));
  orx  g0439(.A(n489), .B(n488), .O(n487));
  andx g0440(.A(n612), .B(po03), .O(n488));
  andx g0441(.A(n490), .B(n614), .O(n489));
  orx  g0442(.A(n53), .B(n618), .O(n490));
  xorx g0443(.A(n493), .B(n74), .O(n491));
  andx g0444(.A(n493), .B(po08), .O(n492));
  orx  g0445(.A(n501), .B(n494), .O(n493));
  invx g0446(.A(n495), .O(n494));
  orx  g0447(.A(n500), .B(n496), .O(n495));
  orx  g0448(.A(n498), .B(n497), .O(n496));
  andx g0449(.A(n621), .B(n102), .O(n497));
  andx g0450(.A(n499), .B(n623), .O(n498));
  orx  g0451(.A(n527), .B(n627), .O(n499));
  xorx g0452(.A(n502), .B(n49), .O(n500));
  andx g0453(.A(n502), .B(n129), .O(n501));
  orx  g0454(.A(n510), .B(n503), .O(n502));
  invx g0455(.A(n504), .O(n503));
  orx  g0456(.A(n509), .B(n505), .O(n504));
  orx  g0457(.A(n507), .B(n506), .O(n505));
  andx g0458(.A(n630), .B(po03), .O(n506));
  andx g0459(.A(n508), .B(n632), .O(n507));
  orx  g0460(.A(n52), .B(n637), .O(n508));
  xorx g0461(.A(n511), .B(n55), .O(n509));
  andx g0462(.A(n511), .B(n78), .O(n510));
  orx  g0463(.A(n519), .B(n512), .O(n511));
  invx g0464(.A(n513), .O(n512));
  orx  g0465(.A(n518), .B(n514), .O(n513));
  orx  g0466(.A(n516), .B(n515), .O(n514));
  andx g0467(.A(n640), .B(n104), .O(n515));
  andx g0468(.A(n643), .B(n517), .O(n516));
  orx  g0469(.A(n53), .B(n642), .O(n517));
  xorx g0470(.A(n520), .B(n57), .O(n518));
  andx g0471(.A(n520), .B(po05), .O(n519));
  orx  g0472(.A(n529), .B(n521), .O(n520));
  invx g0473(.A(n522), .O(n521));
  orx  g0474(.A(n528), .B(n523), .O(n522));
  orx  g0475(.A(n525), .B(n524), .O(n523));
  andx g0476(.A(n645), .B(n104), .O(n524));
  andx g0477(.A(pi07), .B(n526), .O(n525));
  orx  g0478(.A(n527), .B(pi06), .O(n526));
  invx g0479(.A(n104), .O(n527));
  xorx g0480(.A(n530), .B(n72), .O(n528));
  andx g0481(.A(n530), .B(po04), .O(n529));
  orx  g0482(.A(n535), .B(n531), .O(n530));
  invx g0483(.A(n532), .O(n531));
  orx  g0484(.A(n534), .B(n533), .O(n532));
  xorx g0485(.A(n102), .B(n1295), .O(n533));
  xorx g0486(.A(po03), .B(pi06), .O(n534));
  andx g0487(.A(n1294), .B(n102), .O(n535));
  orx  g0488(.A(n647), .B(n537), .O(n536));
  orx  g0489(.A(n539), .B(n538), .O(n537));
  andx g0490(.A(n662), .B(n657), .O(n538));
  andx g0491(.A(n547), .B(n540), .O(n539));
  orx  g0492(.A(n546), .B(n541), .O(n540));
  orx  g0493(.A(n544), .B(n542), .O(n541));
  invx g0494(.A(n543), .O(n542));
  orx  g0495(.A(n664), .B(n73), .O(n543));
  andx g0496(.A(n545), .B(n665), .O(n544));
  orx  g0497(.A(n72), .B(n670), .O(n545));
  xorx g0498(.A(n548), .B(n133), .O(n546));
  orx  g0499(.A(n548), .B(n60), .O(n547));
  andx g0500(.A(n556), .B(n549), .O(n548));
  orx  g0501(.A(n555), .B(n550), .O(n549));
  orx  g0502(.A(n553), .B(n551), .O(n550));
  invx g0503(.A(n552), .O(n551));
  orx  g0504(.A(n673), .B(n73), .O(n552));
  andx g0505(.A(n554), .B(n674), .O(n553));
  orx  g0506(.A(n636), .B(n678), .O(n554));
  xorx g0507(.A(n557), .B(n138), .O(n555));
  orx  g0508(.A(n557), .B(n94), .O(n556));
  andx g0509(.A(n564), .B(n558), .O(n557));
  orx  g0510(.A(n563), .B(n559), .O(n558));
  orx  g0511(.A(n561), .B(n560), .O(n559));
  andx g0512(.A(n682), .B(n124), .O(n560));
  andx g0513(.A(n562), .B(n684), .O(n561));
  orx  g0514(.A(n73), .B(n688), .O(n562));
  xorx g0515(.A(n566), .B(n116), .O(n563));
  invx g0516(.A(n565), .O(n564));
  andx g0517(.A(n566), .B(po13), .O(n565));
  orx  g0518(.A(n574), .B(n567), .O(n566));
  invx g0519(.A(n568), .O(n567));
  orx  g0520(.A(n573), .B(n569), .O(n568));
  orx  g0521(.A(n571), .B(n570), .O(n569));
  andx g0522(.A(n691), .B(n124), .O(n570));
  andx g0523(.A(n572), .B(n693), .O(n571));
  orx  g0524(.A(n72), .B(n697), .O(n572));
  xorx g0525(.A(n575), .B(n71), .O(n573));
  andx g0526(.A(n575), .B(n91), .O(n574));
  orx  g0527(.A(n583), .B(n576), .O(n575));
  invx g0528(.A(n577), .O(n576));
  orx  g0529(.A(n582), .B(n578), .O(n577));
  orx  g0530(.A(n580), .B(n579), .O(n578));
  andx g0531(.A(n700), .B(n122), .O(n579));
  andx g0532(.A(n581), .B(n702), .O(n580));
  orx  g0533(.A(n636), .B(n706), .O(n581));
  xorx g0534(.A(n584), .B(n113), .O(n582));
  andx g0535(.A(n584), .B(n110), .O(n583));
  orx  g0536(.A(n592), .B(n585), .O(n584));
  invx g0537(.A(n586), .O(n585));
  orx  g0538(.A(n591), .B(n587), .O(n586));
  orx  g0539(.A(n589), .B(n588), .O(n587));
  andx g0540(.A(n709), .B(po04), .O(n588));
  andx g0541(.A(n590), .B(n711), .O(n589));
  orx  g0542(.A(n73), .B(n715), .O(n590));
  xorx g0543(.A(n593), .B(n66), .O(n591));
  andx g0544(.A(n593), .B(po10), .O(n592));
  orx  g0545(.A(n601), .B(n594), .O(n593));
  invx g0546(.A(n595), .O(n594));
  orx  g0547(.A(n600), .B(n596), .O(n595));
  orx  g0548(.A(n598), .B(n597), .O(n596));
  andx g0549(.A(n718), .B(n124), .O(n597));
  andx g0550(.A(n599), .B(n720), .O(n598));
  orx  g0551(.A(n72), .B(n724), .O(n599));
  xorx g0552(.A(n602), .B(n62), .O(n600));
  andx g0553(.A(n602), .B(po09), .O(n601));
  orx  g0554(.A(n610), .B(n603), .O(n602));
  invx g0555(.A(n604), .O(n603));
  orx  g0556(.A(n609), .B(n605), .O(n604));
  orx  g0557(.A(n607), .B(n606), .O(n605));
  andx g0558(.A(n727), .B(po04), .O(n606));
  andx g0559(.A(n608), .B(n729), .O(n607));
  orx  g0560(.A(n636), .B(n733), .O(n608));
  xorx g0561(.A(n611), .B(n77), .O(n609));
  andx g0562(.A(n611), .B(n98), .O(n610));
  orx  g0563(.A(n619), .B(n612), .O(n611));
  invx g0564(.A(n613), .O(n612));
  orx  g0565(.A(n618), .B(n614), .O(n613));
  orx  g0566(.A(n616), .B(n615), .O(n614));
  andx g0567(.A(n736), .B(n122), .O(n615));
  andx g0568(.A(n617), .B(n738), .O(n616));
  orx  g0569(.A(n73), .B(n743), .O(n617));
  xorx g0570(.A(n620), .B(n918), .O(n618));
  andx g0571(.A(n620), .B(po07), .O(n619));
  orx  g0572(.A(n628), .B(n621), .O(n620));
  invx g0573(.A(n622), .O(n621));
  orx  g0574(.A(n627), .B(n623), .O(n622));
  orx  g0575(.A(n625), .B(n624), .O(n623));
  andx g0576(.A(n746), .B(po04), .O(n624));
  andx g0577(.A(n749), .B(n626), .O(n625));
  orx  g0578(.A(n72), .B(n748), .O(n626));
  xorx g0579(.A(n629), .B(n54), .O(n627));
  andx g0580(.A(n629), .B(po06), .O(n628));
  orx  g0581(.A(n638), .B(n630), .O(n629));
  invx g0582(.A(n631), .O(n630));
  orx  g0583(.A(n637), .B(n632), .O(n631));
  orx  g0584(.A(n634), .B(n633), .O(n632));
  andx g0585(.A(n1292), .B(n124), .O(n633));
  andx g0586(.A(pi09), .B(n635), .O(n634));
  orx  g0587(.A(n636), .B(pi08), .O(n635));
  invx g0588(.A(n124), .O(n636));
  xorx g0589(.A(n639), .B(n56), .O(n637));
  andx g0590(.A(n639), .B(n101), .O(n638));
  orx  g0591(.A(n644), .B(n640), .O(n639));
  invx g0592(.A(n641), .O(n640));
  orx  g0593(.A(n643), .B(n642), .O(n641));
  xorx g0594(.A(n122), .B(n646), .O(n642));
  xorx g0595(.A(po04), .B(pi08), .O(n643));
  andx g0596(.A(n645), .B(n124), .O(n644));
  invx g0597(.A(n646), .O(n645));
  orx  g0598(.A(pi07), .B(pi06), .O(n646));
  andx g0599(.A(n655), .B(n122), .O(n647));
  orx  g0600(.A(n653), .B(n649), .O(n648));
  orx  g0601(.A(n651), .B(n650), .O(n649));
  andx g0602(.A(n760), .B(n756), .O(n650));
  andx g0603(.A(n652), .B(n656), .O(n651));
  orx  g0604(.A(n663), .B(n61), .O(n652));
  andx g0605(.A(n654), .B(n101), .O(n653));
  invx g0606(.A(n755), .O(n654));
  invx g0607(.A(n656), .O(n655));
  orx  g0608(.A(n662), .B(n657), .O(n656));
  orx  g0609(.A(n660), .B(n658), .O(n657));
  invx g0610(.A(n659), .O(n658));
  orx  g0611(.A(n763), .B(n58), .O(n659));
  andx g0612(.A(n661), .B(n764), .O(n660));
  orx  g0613(.A(n56), .B(n768), .O(n661));
  xorx g0614(.A(n663), .B(n134), .O(n662));
  andx g0615(.A(n671), .B(n664), .O(n663));
  orx  g0616(.A(n670), .B(n665), .O(n664));
  orx  g0617(.A(n668), .B(n666), .O(n665));
  invx g0618(.A(n667), .O(n666));
  orx  g0619(.A(n771), .B(n57), .O(n667));
  andx g0620(.A(n669), .B(n772), .O(n668));
  orx  g0621(.A(n58), .B(n776), .O(n669));
  xorx g0622(.A(n672), .B(po14), .O(n670));
  orx  g0623(.A(n672), .B(n136), .O(n671));
  andx g0624(.A(n679), .B(n673), .O(n672));
  orx  g0625(.A(n678), .B(n674), .O(n673));
  orx  g0626(.A(n676), .B(n675), .O(n674));
  andx g0627(.A(n780), .B(n99), .O(n675));
  andx g0628(.A(n677), .B(n782), .O(n676));
  orx  g0629(.A(n57), .B(n786), .O(n677));
  xorx g0630(.A(n681), .B(n1241), .O(n678));
  invx g0631(.A(n680), .O(n679));
  andx g0632(.A(n681), .B(n106), .O(n680));
  orx  g0633(.A(n689), .B(n682), .O(n681));
  invx g0634(.A(n683), .O(n682));
  orx  g0635(.A(n688), .B(n684), .O(n683));
  orx  g0636(.A(n686), .B(n685), .O(n684));
  andx g0637(.A(n789), .B(po05), .O(n685));
  andx g0638(.A(n687), .B(n791), .O(n686));
  orx  g0639(.A(n56), .B(n795), .O(n687));
  xorx g0640(.A(n690), .B(n70), .O(n688));
  andx g0641(.A(n690), .B(po12), .O(n689));
  orx  g0642(.A(n698), .B(n691), .O(n690));
  invx g0643(.A(n692), .O(n691));
  orx  g0644(.A(n697), .B(n693), .O(n692));
  orx  g0645(.A(n695), .B(n694), .O(n693));
  andx g0646(.A(n798), .B(n101), .O(n694));
  andx g0647(.A(n696), .B(n800), .O(n695));
  orx  g0648(.A(n58), .B(n804), .O(n696));
  xorx g0649(.A(n699), .B(n1168), .O(n697));
  andx g0650(.A(n699), .B(n111), .O(n698));
  orx  g0651(.A(n707), .B(n700), .O(n699));
  invx g0652(.A(n701), .O(n700));
  orx  g0653(.A(n706), .B(n702), .O(n701));
  orx  g0654(.A(n704), .B(n703), .O(n702));
  andx g0655(.A(n807), .B(po05), .O(n703));
  andx g0656(.A(n705), .B(n809), .O(n704));
  orx  g0657(.A(n57), .B(n813), .O(n705));
  xorx g0658(.A(n708), .B(n65), .O(n706));
  andx g0659(.A(n708), .B(n87), .O(n707));
  orx  g0660(.A(n716), .B(n709), .O(n708));
  invx g0661(.A(n710), .O(n709));
  orx  g0662(.A(n715), .B(n711), .O(n710));
  orx  g0663(.A(n713), .B(n712), .O(n711));
  andx g0664(.A(n816), .B(n99), .O(n712));
  andx g0665(.A(n714), .B(n818), .O(n713));
  orx  g0666(.A(n56), .B(n822), .O(n714));
  xorx g0667(.A(n717), .B(n1063), .O(n715));
  andx g0668(.A(n717), .B(n127), .O(n716));
  orx  g0669(.A(n725), .B(n718), .O(n717));
  invx g0670(.A(n719), .O(n718));
  orx  g0671(.A(n724), .B(n720), .O(n719));
  orx  g0672(.A(n722), .B(n721), .O(n720));
  andx g0673(.A(n825), .B(po05), .O(n721));
  andx g0674(.A(n723), .B(n827), .O(n722));
  orx  g0675(.A(n58), .B(n832), .O(n723));
  xorx g0676(.A(n726), .B(n76), .O(n724));
  andx g0677(.A(n726), .B(po08), .O(n725));
  orx  g0678(.A(n734), .B(n727), .O(n726));
  invx g0679(.A(n728), .O(n727));
  orx  g0680(.A(n733), .B(n729), .O(n728));
  orx  g0681(.A(n731), .B(n730), .O(n729));
  andx g0682(.A(n835), .B(n101), .O(n730));
  andx g0683(.A(n838), .B(n732), .O(n731));
  orx  g0684(.A(n57), .B(n837), .O(n732));
  xorx g0685(.A(n735), .B(n48), .O(n733));
  andx g0686(.A(n735), .B(po07), .O(n734));
  orx  g0687(.A(n744), .B(n736), .O(n735));
  invx g0688(.A(n737), .O(n736));
  orx  g0689(.A(n743), .B(n738), .O(n737));
  orx  g0690(.A(n740), .B(n739), .O(n738));
  andx g0691(.A(n840), .B(n101), .O(n739));
  andx g0692(.A(pi11), .B(n741), .O(n740));
  orx  g0693(.A(n56), .B(pi10), .O(n741));
  invx g0694(.A(n101), .O(n742));
  xorx g0695(.A(n745), .B(n831), .O(n743));
  andx g0696(.A(n745), .B(n80), .O(n744));
  orx  g0697(.A(n750), .B(n746), .O(n745));
  invx g0698(.A(n747), .O(n746));
  orx  g0699(.A(n749), .B(n748), .O(n747));
  xorx g0700(.A(n99), .B(n1293), .O(n748));
  xorx g0701(.A(po05), .B(pi10), .O(n749));
  andx g0702(.A(n1292), .B(n99), .O(n750));
  orx  g0703(.A(n842), .B(n752), .O(n751));
  orx  g0704(.A(n754), .B(n753), .O(n752));
  andx g0705(.A(n856), .B(n852), .O(n753));
  andx g0706(.A(n761), .B(n755), .O(n754));
  orx  g0707(.A(n760), .B(n756), .O(n755));
  orx  g0708(.A(n758), .B(n757), .O(n756));
  andx g0709(.A(n858), .B(n80), .O(n757));
  andx g0710(.A(n759), .B(n860), .O(n758));
  orx  g0711(.A(n831), .B(n864), .O(n759));
  xorx g0712(.A(n762), .B(n135), .O(n760));
  orx  g0713(.A(n762), .B(n60), .O(n761));
  andx g0714(.A(n769), .B(n763), .O(n762));
  orx  g0715(.A(n768), .B(n764), .O(n763));
  orx  g0716(.A(n766), .B(n765), .O(n764));
  andx g0717(.A(n867), .B(n78), .O(n765));
  andx g0718(.A(n767), .B(n869), .O(n766));
  orx  g0719(.A(n55), .B(n873), .O(n767));
  xorx g0720(.A(n770), .B(n140), .O(n768));
  orx  g0721(.A(n770), .B(n95), .O(n769));
  andx g0722(.A(n777), .B(n771), .O(n770));
  orx  g0723(.A(n776), .B(n772), .O(n771));
  orx  g0724(.A(n774), .B(n773), .O(n772));
  andx g0725(.A(n876), .B(po06), .O(n773));
  andx g0726(.A(n775), .B(n878), .O(n774));
  orx  g0727(.A(n54), .B(n882), .O(n775));
  xorx g0728(.A(n779), .B(n118), .O(n776));
  invx g0729(.A(n778), .O(n777));
  andx g0730(.A(n779), .B(n107), .O(n778));
  orx  g0731(.A(n787), .B(n780), .O(n779));
  invx g0732(.A(n781), .O(n780));
  orx  g0733(.A(n786), .B(n782), .O(n781));
  orx  g0734(.A(n784), .B(n783), .O(n782));
  andx g0735(.A(n885), .B(n80), .O(n783));
  andx g0736(.A(n785), .B(n887), .O(n784));
  orx  g0737(.A(n54), .B(n891), .O(n785));
  xorx g0738(.A(n788), .B(n69), .O(n786));
  andx g0739(.A(n788), .B(n91), .O(n787));
  orx  g0740(.A(n796), .B(n789), .O(n788));
  invx g0741(.A(n790), .O(n789));
  orx  g0742(.A(n795), .B(n791), .O(n790));
  orx  g0743(.A(n793), .B(n792), .O(n791));
  andx g0744(.A(n894), .B(po06), .O(n792));
  andx g0745(.A(n794), .B(n896), .O(n793));
  orx  g0746(.A(n55), .B(n900), .O(n794));
  xorx g0747(.A(n797), .B(n112), .O(n795));
  andx g0748(.A(n797), .B(n108), .O(n796));
  orx  g0749(.A(n805), .B(n798), .O(n797));
  invx g0750(.A(n799), .O(n798));
  orx  g0751(.A(n804), .B(n800), .O(n799));
  orx  g0752(.A(n802), .B(n801), .O(n800));
  andx g0753(.A(n903), .B(n78), .O(n801));
  andx g0754(.A(n803), .B(n905), .O(n802));
  orx  g0755(.A(n54), .B(n909), .O(n803));
  xorx g0756(.A(n806), .B(n68), .O(n804));
  andx g0757(.A(n806), .B(po10), .O(n805));
  orx  g0758(.A(n814), .B(n807), .O(n806));
  invx g0759(.A(n808), .O(n807));
  orx  g0760(.A(n813), .B(n809), .O(n808));
  orx  g0761(.A(n811), .B(n810), .O(n809));
  andx g0762(.A(n912), .B(po06), .O(n810));
  andx g0763(.A(n812), .B(n914), .O(n811));
  orx  g0764(.A(n55), .B(n919), .O(n812));
  xorx g0765(.A(n815), .B(n64), .O(n813));
  andx g0766(.A(n815), .B(po09), .O(n814));
  orx  g0767(.A(n823), .B(n816), .O(n815));
  invx g0768(.A(n817), .O(n816));
  orx  g0769(.A(n822), .B(n818), .O(n817));
  orx  g0770(.A(n820), .B(n819), .O(n818));
  andx g0771(.A(n922), .B(n80), .O(n819));
  andx g0772(.A(n925), .B(n821), .O(n820));
  orx  g0773(.A(n55), .B(n924), .O(n821));
  xorx g0774(.A(n824), .B(n75), .O(n822));
  andx g0775(.A(n824), .B(n98), .O(n823));
  orx  g0776(.A(n833), .B(n825), .O(n824));
  invx g0777(.A(n826), .O(n825));
  orx  g0778(.A(n832), .B(n827), .O(n826));
  orx  g0779(.A(n829), .B(n828), .O(n827));
  andx g0780(.A(n1290), .B(n80), .O(n828));
  andx g0781(.A(pi13), .B(n830), .O(n829));
  orx  g0782(.A(n54), .B(pi12), .O(n830));
  invx g0783(.A(po06), .O(n831));
  xorx g0784(.A(n930), .B(n834), .O(n832));
  andx g0785(.A(n834), .B(n931), .O(n833));
  orx  g0786(.A(n839), .B(n835), .O(n834));
  invx g0787(.A(n836), .O(n835));
  orx  g0788(.A(n838), .B(n837), .O(n836));
  xorx g0789(.A(n847), .B(n841), .O(n837));
  xorx g0790(.A(n78), .B(pi12), .O(n838));
  andx g0791(.A(n840), .B(n847), .O(n839));
  invx g0792(.A(n841), .O(n840));
  orx  g0793(.A(pi11), .B(pi10), .O(n841));
  andx g0794(.A(n850), .B(n78), .O(n842));
  orx  g0795(.A(n849), .B(n844), .O(n843));
  orx  g0796(.A(n846), .B(n845), .O(n844));
  andx g0797(.A(n939), .B(n934), .O(n845));
  invx g0798(.A(n847), .O(n846));
  orx  g0799(.A(n848), .B(n850), .O(n847));
  andx g0800(.A(n857), .B(n135), .O(n848));
  andx g0801(.A(n932), .B(n128), .O(n849));
  invx g0802(.A(n851), .O(n850));
  orx  g0803(.A(n856), .B(n852), .O(n851));
  orx  g0804(.A(n854), .B(n853), .O(n852));
  andx g0805(.A(n942), .B(n129), .O(n853));
  andx g0806(.A(n855), .B(n944), .O(n854));
  orx  g0807(.A(n49), .B(n949), .O(n855));
  xorx g0808(.A(n857), .B(n59), .O(n856));
  orx  g0809(.A(n865), .B(n858), .O(n857));
  invx g0810(.A(n859), .O(n858));
  orx  g0811(.A(n864), .B(n860), .O(n859));
  orx  g0812(.A(n862), .B(n861), .O(n860));
  andx g0813(.A(n952), .B(po07), .O(n861));
  andx g0814(.A(n863), .B(n954), .O(n862));
  orx  g0815(.A(n918), .B(n958), .O(n863));
  xorx g0816(.A(n866), .B(n94), .O(n864));
  andx g0817(.A(n866), .B(n137), .O(n865));
  orx  g0818(.A(n874), .B(n867), .O(n866));
  invx g0819(.A(n868), .O(n867));
  orx  g0820(.A(n873), .B(n869), .O(n868));
  orx  g0821(.A(n871), .B(n870), .O(n869));
  andx g0822(.A(n961), .B(po07), .O(n870));
  andx g0823(.A(n872), .B(n963), .O(n871));
  orx  g0824(.A(n48), .B(n967), .O(n872));
  xorx g0825(.A(n875), .B(n117), .O(n873));
  andx g0826(.A(n875), .B(po13), .O(n874));
  orx  g0827(.A(n883), .B(n876), .O(n875));
  invx g0828(.A(n877), .O(n876));
  orx  g0829(.A(n882), .B(n878), .O(n877));
  orx  g0830(.A(n880), .B(n879), .O(n878));
  andx g0831(.A(n970), .B(n128), .O(n879));
  andx g0832(.A(n881), .B(n972), .O(n880));
  orx  g0833(.A(n49), .B(n976), .O(n881));
  xorx g0834(.A(n884), .B(n88), .O(n882));
  andx g0835(.A(n884), .B(po12), .O(n883));
  orx  g0836(.A(n892), .B(n885), .O(n884));
  invx g0837(.A(n886), .O(n885));
  orx  g0838(.A(n891), .B(n887), .O(n886));
  orx  g0839(.A(n889), .B(n888), .O(n887));
  andx g0840(.A(n979), .B(n129), .O(n888));
  andx g0841(.A(n890), .B(n981), .O(n889));
  orx  g0842(.A(n49), .B(n985), .O(n890));
  xorx g0843(.A(n893), .B(n114), .O(n891));
  andx g0844(.A(n893), .B(n109), .O(n892));
  orx  g0845(.A(n901), .B(n894), .O(n893));
  invx g0846(.A(n895), .O(n894));
  orx  g0847(.A(n900), .B(n896), .O(n895));
  orx  g0848(.A(n898), .B(n897), .O(n896));
  andx g0849(.A(n988), .B(po07), .O(n897));
  andx g0850(.A(n899), .B(n990), .O(n898));
  orx  g0851(.A(n48), .B(n994), .O(n899));
  xorx g0852(.A(n902), .B(n67), .O(n900));
  andx g0853(.A(n902), .B(n87), .O(n901));
  orx  g0854(.A(n910), .B(n903), .O(n902));
  invx g0855(.A(n904), .O(n903));
  orx  g0856(.A(n909), .B(n905), .O(n904));
  orx  g0857(.A(n907), .B(n906), .O(n905));
  andx g0858(.A(n997), .B(n129), .O(n906));
  andx g0859(.A(n1000), .B(n908), .O(n907));
  orx  g0860(.A(n49), .B(n999), .O(n908));
  xorx g0861(.A(n911), .B(n63), .O(n909));
  andx g0862(.A(n911), .B(n127), .O(n910));
  orx  g0863(.A(n920), .B(n912), .O(n911));
  invx g0864(.A(n913), .O(n912));
  orx  g0865(.A(n919), .B(n914), .O(n913));
  orx  g0866(.A(n916), .B(n915), .O(n914));
  andx g0867(.A(n1002), .B(n128), .O(n915));
  andx g0868(.A(pi15), .B(n917), .O(n916));
  orx  g0869(.A(n918), .B(pi14), .O(n917));
  invx g0870(.A(po07), .O(n918));
  xorx g0871(.A(n921), .B(n74), .O(n919));
  andx g0872(.A(n921), .B(po08), .O(n920));
  orx  g0873(.A(n926), .B(n922), .O(n921));
  invx g0874(.A(n923), .O(n922));
  orx  g0875(.A(n925), .B(n924), .O(n923));
  xorx g0876(.A(n128), .B(n1291), .O(n924));
  xorx g0877(.A(n129), .B(pi14), .O(n925));
  andx g0878(.A(n1290), .B(n129), .O(n926));
  orx  g0879(.A(n1004), .B(n928), .O(n927));
  orx  g0880(.A(n930), .B(n929), .O(n928));
  andx g0881(.A(n1019), .B(n1014), .O(n929));
  invx g0882(.A(n931), .O(n930));
  orx  g0883(.A(n940), .B(n932), .O(n931));
  invx g0884(.A(n933), .O(n932));
  orx  g0885(.A(n939), .B(n934), .O(n933));
  orx  g0886(.A(n937), .B(n935), .O(n934));
  invx g0887(.A(n936), .O(n935));
  orx  g0888(.A(n1021), .B(n77), .O(n936));
  andx g0889(.A(n938), .B(n1022), .O(n937));
  orx  g0890(.A(n74), .B(n1027), .O(n938));
  xorx g0891(.A(n941), .B(n59), .O(n939));
  andx g0892(.A(n941), .B(po15), .O(n940));
  orx  g0893(.A(n950), .B(n942), .O(n941));
  invx g0894(.A(n943), .O(n942));
  orx  g0895(.A(n949), .B(n944), .O(n943));
  orx  g0896(.A(n947), .B(n945), .O(n944));
  invx g0897(.A(n946), .O(n945));
  orx  g0898(.A(n1030), .B(n76), .O(n946));
  andx g0899(.A(n948), .B(n1031), .O(n947));
  orx  g0900(.A(n77), .B(n1035), .O(n948));
  xorx g0901(.A(n951), .B(n1266), .O(n949));
  andx g0902(.A(n951), .B(n138), .O(n950));
  orx  g0903(.A(n959), .B(n952), .O(n951));
  invx g0904(.A(n953), .O(n952));
  orx  g0905(.A(n958), .B(n954), .O(n953));
  orx  g0906(.A(n956), .B(n955), .O(n954));
  andx g0907(.A(n1039), .B(n98), .O(n955));
  andx g0908(.A(n957), .B(n1041), .O(n956));
  orx  g0909(.A(n76), .B(n1045), .O(n957));
  xorx g0910(.A(n960), .B(n116), .O(n958));
  andx g0911(.A(n960), .B(n106), .O(n959));
  orx  g0912(.A(n968), .B(n961), .O(n960));
  invx g0913(.A(n962), .O(n961));
  orx  g0914(.A(n967), .B(n963), .O(n962));
  orx  g0915(.A(n965), .B(n964), .O(n963));
  andx g0916(.A(n1048), .B(po08), .O(n964));
  andx g0917(.A(n966), .B(n1050), .O(n965));
  orx  g0918(.A(n75), .B(n1054), .O(n966));
  xorx g0919(.A(n969), .B(n71), .O(n967));
  andx g0920(.A(n969), .B(n91), .O(n968));
  orx  g0921(.A(n977), .B(n970), .O(n969));
  invx g0922(.A(n971), .O(n970));
  orx  g0923(.A(n976), .B(n972), .O(n971));
  orx  g0924(.A(n974), .B(n973), .O(n972));
  andx g0925(.A(n1057), .B(n98), .O(n973));
  andx g0926(.A(n975), .B(n1059), .O(n974));
  orx  g0927(.A(n74), .B(n1064), .O(n975));
  xorx g0928(.A(n978), .B(n113), .O(n976));
  andx g0929(.A(n978), .B(n110), .O(n977));
  orx  g0930(.A(n986), .B(n979), .O(n978));
  invx g0931(.A(n980), .O(n979));
  orx  g0932(.A(n985), .B(n981), .O(n980));
  orx  g0933(.A(n983), .B(n982), .O(n981));
  andx g0934(.A(n1067), .B(po08), .O(n982));
  andx g0935(.A(n1070), .B(n984), .O(n983));
  orx  g0936(.A(n77), .B(n1069), .O(n984));
  xorx g0937(.A(n987), .B(n66), .O(n985));
  andx g0938(.A(n987), .B(po10), .O(n986));
  orx  g0939(.A(n995), .B(n988), .O(n987));
  invx g0940(.A(n989), .O(n988));
  orx  g0941(.A(n994), .B(n990), .O(n989));
  orx  g0942(.A(n992), .B(n991), .O(n990));
  andx g0943(.A(n1288), .B(n98), .O(n991));
  andx g0944(.A(pi17), .B(n993), .O(n992));
  orx  g0945(.A(n76), .B(pi16), .O(n993));
  xorx g0946(.A(n996), .B(n62), .O(n994));
  andx g0947(.A(n996), .B(po09), .O(n995));
  orx  g0948(.A(n1001), .B(n997), .O(n996));
  invx g0949(.A(n998), .O(n997));
  orx  g0950(.A(n1000), .B(n999), .O(n998));
  xorx g0951(.A(n1006), .B(n1003), .O(n999));
  xorx g0952(.A(n1006), .B(pi16), .O(n1000));
  andx g0953(.A(n1002), .B(po08), .O(n1001));
  invx g0954(.A(n1003), .O(n1002));
  orx  g0955(.A(pi15), .B(pi14), .O(n1003));
  invx g0956(.A(n1005), .O(n1004));
  orx  g0957(.A(n1013), .B(n75), .O(n1005));
  orx  g0958(.A(n1011), .B(n1007), .O(n1006));
  orx  g0959(.A(n1009), .B(n1008), .O(n1007));
  andx g0960(.A(n1082), .B(n1077), .O(n1008));
  andx g0961(.A(n1010), .B(n1013), .O(n1009));
  orx  g0962(.A(n1020), .B(n61), .O(n1010));
  andx g0963(.A(n1012), .B(n127), .O(n1011));
  invx g0964(.A(n1076), .O(n1012));
  orx  g0965(.A(n1019), .B(n1014), .O(n1013));
  orx  g0966(.A(n1017), .B(n1015), .O(n1014));
  invx g0967(.A(n1016), .O(n1015));
  orx  g0968(.A(n1085), .B(n64), .O(n1016));
  andx g0969(.A(n1018), .B(n1086), .O(n1017));
  orx  g0970(.A(n62), .B(n1091), .O(n1018));
  xorx g0971(.A(n1020), .B(po15), .O(n1019));
  andx g0972(.A(n1028), .B(n1021), .O(n1020));
  orx  g0973(.A(n1027), .B(n1022), .O(n1021));
  orx  g0974(.A(n1025), .B(n1023), .O(n1022));
  invx g0975(.A(n1024), .O(n1023));
  orx  g0976(.A(n1094), .B(n63), .O(n1024));
  andx g0977(.A(n1026), .B(n1095), .O(n1025));
  orx  g0978(.A(n1063), .B(n1099), .O(n1026));
  xorx g0979(.A(n1029), .B(n137), .O(n1027));
  orx  g0980(.A(n1029), .B(n94), .O(n1028));
  andx g0981(.A(n1036), .B(n1030), .O(n1029));
  orx  g0982(.A(n1035), .B(n1031), .O(n1030));
  orx  g0983(.A(n1033), .B(n1032), .O(n1031));
  andx g0984(.A(n1103), .B(po09), .O(n1032));
  andx g0985(.A(n1034), .B(n1105), .O(n1033));
  orx  g0986(.A(n64), .B(n1109), .O(n1034));
  xorx g0987(.A(n1038), .B(n1241), .O(n1035));
  invx g0988(.A(n1037), .O(n1036));
  andx g0989(.A(n1038), .B(n107), .O(n1037));
  orx  g0990(.A(n1046), .B(n1039), .O(n1038));
  invx g0991(.A(n1040), .O(n1039));
  orx  g0992(.A(n1045), .B(n1041), .O(n1040));
  orx  g0993(.A(n1043), .B(n1042), .O(n1041));
  andx g0994(.A(n1112), .B(n127), .O(n1042));
  andx g0995(.A(n1044), .B(n1114), .O(n1043));
  orx  g0996(.A(n63), .B(n1118), .O(n1044));
  xorx g0997(.A(n1047), .B(n70), .O(n1045));
  andx g0998(.A(n1047), .B(po12), .O(n1046));
  orx  g0999(.A(n1055), .B(n1048), .O(n1047));
  invx g1000(.A(n1049), .O(n1048));
  orx  g1001(.A(n1054), .B(n1050), .O(n1049));
  orx  g1002(.A(n1052), .B(n1051), .O(n1050));
  andx g1003(.A(n1121), .B(po09), .O(n1051));
  andx g1004(.A(n1124), .B(n1053), .O(n1052));
  orx  g1005(.A(n62), .B(n1123), .O(n1053));
  xorx g1006(.A(n1056), .B(n1168), .O(n1054));
  andx g1007(.A(n1056), .B(n110), .O(n1055));
  orx  g1008(.A(n1065), .B(n1057), .O(n1056));
  invx g1009(.A(n1058), .O(n1057));
  orx  g1010(.A(n1064), .B(n1059), .O(n1058));
  orx  g1011(.A(n1061), .B(n1060), .O(n1059));
  andx g1012(.A(n1126), .B(n127), .O(n1060));
  andx g1013(.A(pi19), .B(n1062), .O(n1061));
  orx  g1014(.A(n1063), .B(pi18), .O(n1062));
  invx g1015(.A(n125), .O(n1063));
  xorx g1016(.A(n1066), .B(n65), .O(n1064));
  andx g1017(.A(n1066), .B(n87), .O(n1065));
  orx  g1018(.A(n1071), .B(n1067), .O(n1066));
  invx g1019(.A(n1068), .O(n1067));
  orx  g1020(.A(n1070), .B(n1069), .O(n1068));
  xorx g1021(.A(n125), .B(n1289), .O(n1069));
  xorx g1022(.A(n125), .B(pi18), .O(n1070));
  andx g1023(.A(n1288), .B(po09), .O(n1071));
  orx  g1024(.A(n1128), .B(n1073), .O(n1072));
  orx  g1025(.A(n1075), .B(n1074), .O(n1073));
  andx g1026(.A(n1143), .B(n1139), .O(n1074));
  andx g1027(.A(n1083), .B(n1076), .O(n1075));
  orx  g1028(.A(n1082), .B(n1077), .O(n1076));
  orx  g1029(.A(n1080), .B(n1078), .O(n1077));
  invx g1030(.A(n1079), .O(n1078));
  orx  g1031(.A(n1145), .B(n67), .O(n1079));
  andx g1032(.A(n1081), .B(n1146), .O(n1080));
  orx  g1033(.A(n65), .B(n1150), .O(n1081));
  xorx g1034(.A(n1084), .B(n133), .O(n1082));
  orx  g1035(.A(n1084), .B(n60), .O(n1083));
  andx g1036(.A(n1092), .B(n1085), .O(n1084));
  orx  g1037(.A(n1091), .B(n1086), .O(n1085));
  orx  g1038(.A(n1089), .B(n1087), .O(n1086));
  invx g1039(.A(n1088), .O(n1087));
  orx  g1040(.A(n1153), .B(n66), .O(n1088));
  andx g1041(.A(n1090), .B(n1154), .O(n1089));
  orx  g1042(.A(n68), .B(n1158), .O(n1090));
  xorx g1043(.A(n1093), .B(n138), .O(n1091));
  orx  g1044(.A(n1093), .B(n136), .O(n1092));
  andx g1045(.A(n1100), .B(n1094), .O(n1093));
  orx  g1046(.A(n1099), .B(n1095), .O(n1094));
  orx  g1047(.A(n1097), .B(n1096), .O(n1095));
  andx g1048(.A(n1162), .B(po10), .O(n1096));
  andx g1049(.A(n1098), .B(n1164), .O(n1097));
  orx  g1050(.A(n67), .B(n1169), .O(n1098));
  xorx g1051(.A(n1102), .B(n118), .O(n1099));
  invx g1052(.A(n1101), .O(n1100));
  andx g1053(.A(n1102), .B(po13), .O(n1101));
  orx  g1054(.A(n1110), .B(n1103), .O(n1102));
  invx g1055(.A(n1104), .O(n1103));
  orx  g1056(.A(n1109), .B(n1105), .O(n1104));
  orx  g1057(.A(n1107), .B(n1106), .O(n1105));
  andx g1058(.A(n1172), .B(n87), .O(n1106));
  andx g1059(.A(n1175), .B(n1108), .O(n1107));
  orx  g1060(.A(n66), .B(n1174), .O(n1108));
  xorx g1061(.A(n1111), .B(n69), .O(n1109));
  andx g1062(.A(n1111), .B(n91), .O(n1110));
  orx  g1063(.A(n1119), .B(n1112), .O(n1111));
  invx g1064(.A(n1113), .O(n1112));
  orx  g1065(.A(n1118), .B(n1114), .O(n1113));
  orx  g1066(.A(n1116), .B(n1115), .O(n1114));
  andx g1067(.A(n1286), .B(po10), .O(n1115));
  andx g1068(.A(pi21), .B(n1117), .O(n1116));
  orx  g1069(.A(n65), .B(pi20), .O(n1117));
  xorx g1070(.A(n1120), .B(n112), .O(n1118));
  andx g1071(.A(n1120), .B(n108), .O(n1119));
  orx  g1072(.A(n1125), .B(n1121), .O(n1120));
  invx g1073(.A(n1122), .O(n1121));
  orx  g1074(.A(n1124), .B(n1123), .O(n1122));
  xorx g1075(.A(n85), .B(n1127), .O(n1123));
  xorx g1076(.A(n85), .B(pi20), .O(n1124));
  andx g1077(.A(n1126), .B(n87), .O(n1125));
  invx g1078(.A(n1127), .O(n1126));
  orx  g1079(.A(pi19), .B(pi18), .O(n1127));
  andx g1080(.A(n1137), .B(po10), .O(n1128));
  orx  g1081(.A(n1135), .B(n1130), .O(n1129));
  orx  g1082(.A(n1133), .B(n1131), .O(n1130));
  andx g1083(.A(n1132), .B(n1190), .O(n1131));
  andx g1084(.A(n1183), .B(n133), .O(n1132));
  andx g1085(.A(n1134), .B(n1138), .O(n1133));
  orx  g1086(.A(n1144), .B(n61), .O(n1134));
  andx g1087(.A(n1136), .B(n109), .O(n1135));
  invx g1088(.A(n1182), .O(n1136));
  invx g1089(.A(n1138), .O(n1137));
  orx  g1090(.A(n1143), .B(n1139), .O(n1138));
  orx  g1091(.A(n1141), .B(n1140), .O(n1139));
  andx g1092(.A(n1191), .B(n110), .O(n1140));
  andx g1093(.A(n1142), .B(n1193), .O(n1141));
  orx  g1094(.A(n112), .B(n1197), .O(n1142));
  xorx g1095(.A(n1144), .B(n134), .O(n1143));
  andx g1096(.A(n1151), .B(n1145), .O(n1144));
  orx  g1097(.A(n1150), .B(n1146), .O(n1145));
  orx  g1098(.A(n1148), .B(n1147), .O(n1146));
  andx g1099(.A(n1200), .B(n109), .O(n1147));
  andx g1100(.A(n1149), .B(n1202), .O(n1148));
  orx  g1101(.A(n114), .B(n1206), .O(n1149));
  xorx g1102(.A(n1152), .B(po14), .O(n1150));
  orx  g1103(.A(n1152), .B(n95), .O(n1151));
  andx g1104(.A(n1159), .B(n1153), .O(n1152));
  orx  g1105(.A(n1158), .B(n1154), .O(n1153));
  orx  g1106(.A(n1156), .B(n1155), .O(n1154));
  andx g1107(.A(n1209), .B(n108), .O(n1155));
  andx g1108(.A(n1212), .B(n1157), .O(n1156));
  orx  g1109(.A(n113), .B(n1211), .O(n1157));
  xorx g1110(.A(n1161), .B(n117), .O(n1158));
  invx g1111(.A(n1160), .O(n1159));
  andx g1112(.A(n1161), .B(n106), .O(n1160));
  orx  g1113(.A(n1170), .B(n1162), .O(n1161));
  invx g1114(.A(n1163), .O(n1162));
  orx  g1115(.A(n1169), .B(n1164), .O(n1163));
  orx  g1116(.A(n1166), .B(n1165), .O(n1164));
  andx g1117(.A(n1214), .B(n109), .O(n1165));
  andx g1118(.A(pi23), .B(n1167), .O(n1166));
  orx  g1119(.A(n114), .B(pi22), .O(n1167));
  invx g1120(.A(n110), .O(n1168));
  xorx g1121(.A(n1171), .B(n1218), .O(n1169));
  andx g1122(.A(n1171), .B(po12), .O(n1170));
  orx  g1123(.A(n1176), .B(n1172), .O(n1171));
  invx g1124(.A(n1173), .O(n1172));
  orx  g1125(.A(n1175), .B(n1174), .O(n1173));
  xorx g1126(.A(n108), .B(n1287), .O(n1174));
  xorx g1127(.A(n109), .B(pi22), .O(n1175));
  andx g1128(.A(n1286), .B(n110), .O(n1176));
  orx  g1129(.A(n1216), .B(n1178), .O(po11));
  orx  g1130(.A(n1181), .B(n1179), .O(n1178));
  andx g1131(.A(n1180), .B(n1234), .O(n1179));
  andx g1132(.A(n1229), .B(n134), .O(n1180));
  andx g1133(.A(n1188), .B(n1182), .O(n1181));
  orx  g1134(.A(n1187), .B(n1183), .O(n1182));
  orx  g1135(.A(n1185), .B(n1184), .O(n1183));
  andx g1136(.A(n1235), .B(n91), .O(n1184));
  andx g1137(.A(n1186), .B(n1237), .O(n1185));
  orx  g1138(.A(n71), .B(n1242), .O(n1186));
  xorx g1139(.A(n1189), .B(n135), .O(n1187));
  orx  g1140(.A(n1189), .B(n60), .O(n1188));
  invx g1141(.A(n1190), .O(n1189));
  orx  g1142(.A(n1198), .B(n1191), .O(n1190));
  invx g1143(.A(n1192), .O(n1191));
  orx  g1144(.A(n1197), .B(n1193), .O(n1192));
  orx  g1145(.A(n1195), .B(n1194), .O(n1193));
  andx g1146(.A(n1245), .B(po12), .O(n1194));
  andx g1147(.A(n1248), .B(n1196), .O(n1195));
  orx  g1148(.A(n71), .B(n1247), .O(n1196));
  xorx g1149(.A(n1199), .B(n95), .O(n1197));
  andx g1150(.A(n1199), .B(po14), .O(n1198));
  orx  g1151(.A(n1207), .B(n1200), .O(n1199));
  invx g1152(.A(n1201), .O(n1200));
  orx  g1153(.A(n1206), .B(n1202), .O(n1201));
  orx  g1154(.A(n1204), .B(n1203), .O(n1202));
  andx g1155(.A(n1284), .B(n91), .O(n1203));
  andx g1156(.A(pi25), .B(n1205), .O(n1204));
  orx  g1157(.A(n70), .B(pi24), .O(n1205));
  xorx g1158(.A(n1208), .B(n116), .O(n1206));
  andx g1159(.A(n1208), .B(n107), .O(n1207));
  orx  g1160(.A(n1213), .B(n1209), .O(n1208));
  invx g1161(.A(n1210), .O(n1209));
  orx  g1162(.A(n1212), .B(n1211), .O(n1210));
  xorx g1163(.A(n89), .B(n1215), .O(n1211));
  xorx g1164(.A(n89), .B(pi24), .O(n1212));
  andx g1165(.A(n1214), .B(po12), .O(n1213));
  invx g1166(.A(n1215), .O(n1214));
  orx  g1167(.A(pi23), .B(pi22), .O(n1215));
  invx g1168(.A(n1217), .O(n1216));
  orx  g1169(.A(n1228), .B(n69), .O(n1217));
  invx g1170(.A(n89), .O(n1218));
  orx  g1171(.A(n1226), .B(n1220), .O(n1219));
  orx  g1172(.A(n1223), .B(n1221), .O(n1220));
  andx g1173(.A(n1222), .B(n1261), .O(n1221));
  andx g1174(.A(n1270), .B(n135), .O(n1222));
  andx g1175(.A(n1224), .B(n1228), .O(n1223));
  orx  g1176(.A(n1225), .B(n61), .O(n1224));
  invx g1177(.A(n1234), .O(n1225));
  invx g1178(.A(n1227), .O(n1226));
  orx  g1179(.A(n1260), .B(n117), .O(n1227));
  orx  g1180(.A(n1233), .B(n1229), .O(n1228));
  orx  g1181(.A(n1231), .B(n1230), .O(n1229));
  andx g1182(.A(n1271), .B(po13), .O(n1230));
  andx g1183(.A(n1274), .B(n1232), .O(n1231));
  orx  g1184(.A(n116), .B(n1273), .O(n1232));
  xorx g1185(.A(n1234), .B(n59), .O(n1233));
  orx  g1186(.A(n1243), .B(n1235), .O(n1234));
  invx g1187(.A(n1236), .O(n1235));
  orx  g1188(.A(n1242), .B(n1237), .O(n1236));
  orx  g1189(.A(n1239), .B(n1238), .O(n1237));
  andx g1190(.A(n1282), .B(n106), .O(n1238));
  andx g1191(.A(pi27), .B(n1240), .O(n1239));
  orx  g1192(.A(n1241), .B(pi26), .O(n1240));
  invx g1193(.A(n107), .O(n1241));
  xorx g1194(.A(n1244), .B(n94), .O(n1242));
  andx g1195(.A(n1244), .B(n140), .O(n1243));
  orx  g1196(.A(n1249), .B(n1245), .O(n1244));
  invx g1197(.A(n1246), .O(n1245));
  orx  g1198(.A(n1248), .B(n1247), .O(n1246));
  xorx g1199(.A(po13), .B(n1285), .O(n1247));
  xorx g1200(.A(n106), .B(pi26), .O(n1248));
  andx g1201(.A(n1284), .B(n107), .O(n1249));
  orx  g1202(.A(n1254), .B(n1251), .O(n1250));
  orx  g1203(.A(n1253), .B(n1252), .O(n1251));
  andx g1204(.A(n1280), .B(n137), .O(n1252));
  andx g1205(.A(n1269), .B(n1260), .O(n1253));
  orx  g1206(.A(n1258), .B(n1255), .O(n1254));
  invx g1207(.A(n1256), .O(n1255));
  orx  g1208(.A(n1257), .B(n60), .O(n1256));
  orx  g1209(.A(n1281), .B(pi30), .O(n1257));
  andx g1210(.A(n1260), .B(n60), .O(n1258));
  invx g1211(.A(n133), .O(n1259));
  orx  g1212(.A(n1267), .B(n1261), .O(n1260));
  orx  g1213(.A(n1264), .B(n1262), .O(n1261));
  invx g1214(.A(n1263), .O(n1262));
  orx  g1215(.A(n1281), .B(n94), .O(n1263));
  andx g1216(.A(pi29), .B(n1265), .O(n1264));
  orx  g1217(.A(n1266), .B(pi28), .O(n1265));
  invx g1218(.A(n138), .O(n1266));
  xorx g1219(.A(n1269), .B(po15), .O(n1267));
  orx  g1220(.A(pi31), .B(pi30), .O(n1268));
  invx g1221(.A(n1270), .O(n1269));
  orx  g1222(.A(n1275), .B(n1271), .O(n1270));
  invx g1223(.A(n1272), .O(n1271));
  orx  g1224(.A(n1274), .B(n1273), .O(n1272));
  xorx g1225(.A(n140), .B(n1283), .O(n1273));
  xorx g1226(.A(n137), .B(pi28), .O(n1274));
  andx g1227(.A(n1282), .B(n138), .O(n1275));
  orx  g1228(.A(n1278), .B(n1277), .O(n1276));
  andx g1229(.A(pi31), .B(pi30), .O(n1277));
  andx g1230(.A(n1281), .B(n1279), .O(n1278));
  invx g1231(.A(n1280), .O(n1279));
  andx g1232(.A(n1281), .B(pi30), .O(n1280));
  orx  g1233(.A(pi28), .B(pi29), .O(n1281));
  invx g1234(.A(n1283), .O(n1282));
  orx  g1235(.A(pi27), .B(pi26), .O(n1283));
  invx g1236(.A(n1285), .O(n1284));
  orx  g1237(.A(pi25), .B(pi24), .O(n1285));
  invx g1238(.A(n1287), .O(n1286));
  orx  g1239(.A(pi21), .B(pi20), .O(n1287));
  invx g1240(.A(n1289), .O(n1288));
  orx  g1241(.A(pi17), .B(pi16), .O(n1289));
  invx g1242(.A(n1291), .O(n1290));
  orx  g1243(.A(pi13), .B(pi12), .O(n1291));
  invx g1244(.A(n1293), .O(n1292));
  orx  g1245(.A(pi09), .B(pi08), .O(n1293));
  invx g1246(.A(n1295), .O(n1294));
  orx  g1247(.A(pi05), .B(pi04), .O(n1295));
endmodule


