// Benchmark "unsigned_mult" written by ABC on Fri Feb  7 13:47:09 2014

module unsigned_mult ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n33, n34, n36, n37, n38, n40, n41, n42, n43, n44, n46, n47, n48, n49,
    n50, n51, n52, n54, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65,
    n67, n68, n69, n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n81,
    n83, n84, n85, n86, n87, n89, n90, n91, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
    n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723;
  andx g000(.A(n33), .B(n245), .O(po09));
  orx  g001(.A(n34), .B(n314), .O(n33));
  andx g002(.A(n460), .B(n381), .O(n34));
  orx  g003(.A(n37), .B(n36), .O(po08));
  andx g004(.A(n461), .B(n381), .O(n36));
  andx g005(.A(n38), .B(n460), .O(n37));
  invx g006(.A(n381), .O(n38));
  orx  g007(.A(n41), .B(n40), .O(po07));
  andx g008(.A(n451), .B(n43), .O(n40));
  invx g009(.A(n42), .O(n41));
  orx  g010(.A(n43), .B(n451), .O(n42));
  orx  g011(.A(n382), .B(n44), .O(n43));
  invx g012(.A(n384), .O(n44));
  andx g013(.A(n47), .B(n46), .O(po06));
  orx  g014(.A(n444), .B(n49), .O(n46));
  orx  g015(.A(n48), .B(n443), .O(n47));
  invx g016(.A(n49), .O(n48));
  orx  g017(.A(n50), .B(n386), .O(n49));
  andx g018(.A(n52), .B(n51), .O(n50));
  orx  g019(.A(n415), .B(n525), .O(n51));
  invx g020(.A(n389), .O(n52));
  orx  g021(.A(n55), .B(n54), .O(po05));
  andx g022(.A(n434), .B(n57), .O(n54));
  invx g023(.A(n56), .O(n55));
  orx  g024(.A(n57), .B(n434), .O(n56));
  orx  g025(.A(n390), .B(n58), .O(n57));
  invx g026(.A(n392), .O(n58));
  orx  g027(.A(n61), .B(n60), .O(po04));
  andx g028(.A(n427), .B(n63), .O(n60));
  invx g029(.A(n62), .O(n61));
  orx  g030(.A(n63), .B(n427), .O(n62));
  orx  g031(.A(n64), .B(n394), .O(n63));
  andx g032(.A(n398), .B(n65), .O(n64));
  orx  g033(.A(n415), .B(n631), .O(n65));
  orx  g034(.A(n69), .B(n67), .O(po03));
  invx g035(.A(n68), .O(n67));
  orx  g036(.A(n417), .B(n70), .O(n68));
  andx g037(.A(n70), .B(n417), .O(n69));
  andx g038(.A(n399), .B(n71), .O(n70));
  invx g039(.A(n401), .O(n71));
  orx  g040(.A(n81), .B(n73), .O(po02));
  orx  g041(.A(n75), .B(n74), .O(n73));
  andx g042(.A(n77), .B(n406), .O(n74));
  andx g043(.A(n78), .B(n76), .O(n75));
  invx g044(.A(n77), .O(n76));
  andx g045(.A(n412), .B(n411), .O(n77));
  andx g046(.A(n80), .B(n79), .O(n78));
  orx  g047(.A(n411), .B(n412), .O(n79));
  invx g048(.A(n406), .O(n80));
  andx g049(.A(n405), .B(n413), .O(n81));
  orx  g050(.A(n84), .B(n83), .O(po01));
  andx g051(.A(n86), .B(n87), .O(n83));
  invx g052(.A(n85), .O(n84));
  orx  g053(.A(n87), .B(n86), .O(n85));
  andx g054(.A(pi00), .B(pi03), .O(n86));
  orx  g055(.A(n415), .B(n721), .O(n87));
  orx  g056(.A(n103), .B(n89), .O(po15));
  orx  g057(.A(n91), .B(n90), .O(n89));
  andx g058(.A(n96), .B(n98), .O(n90));
  invx g059(.A(n95), .O(n91));
  orx  g060(.A(n97), .B(n93), .O(po14));
  andx g061(.A(n94), .B(n99), .O(n93));
  andx g062(.A(n96), .B(n95), .O(n94));
  orx  g063(.A(n102), .B(n110), .O(n95));
  invx g064(.A(n101), .O(n96));
  andx g065(.A(n101), .B(n98), .O(n97));
  invx g066(.A(n99), .O(n98));
  andx g067(.A(n100), .B(n120), .O(n99));
  orx  g068(.A(n121), .B(n116), .O(n100));
  andx g069(.A(n110), .B(n102), .O(n101));
  orx  g070(.A(n104), .B(n103), .O(n102));
  andx g071(.A(pi02), .B(n107), .O(n103));
  andx g072(.A(n106), .B(n105), .O(n104));
  orx  g073(.A(n303), .B(n504), .O(n105));
  invx g074(.A(n107), .O(n106));
  orx  g075(.A(n108), .B(n133), .O(n107));
  andx g076(.A(n109), .B(pi15), .O(n108));
  andx g077(.A(pi13), .B(n131), .O(n109));
  orx  g078(.A(n126), .B(n111), .O(n110));
  invx g079(.A(n139), .O(n111));
  andx g080(.A(n114), .B(n113), .O(po13));
  orx  g081(.A(n116), .B(n118), .O(n113));
  invx g082(.A(n115), .O(n114));
  andx g083(.A(n118), .B(n116), .O(n115));
  andx g084(.A(n117), .B(n147), .O(n116));
  orx  g085(.A(n152), .B(n145), .O(n117));
  orx  g086(.A(n121), .B(n119), .O(n118));
  invx g087(.A(n120), .O(n119));
  orx  g088(.A(n122), .B(n156), .O(n120));
  andx g089(.A(n156), .B(n122), .O(n121));
  andx g090(.A(n125), .B(n123), .O(n122));
  invx g091(.A(n124), .O(n123));
  andx g092(.A(n126), .B(n139), .O(n124));
  orx  g093(.A(n139), .B(n126), .O(n125));
  orx  g094(.A(n129), .B(n127), .O(n126));
  invx g095(.A(n128), .O(n127));
  orx  g096(.A(n130), .B(n138), .O(n128));
  andx g097(.A(n138), .B(n130), .O(n129));
  andx g098(.A(n132), .B(n131), .O(n130));
  orx  g099(.A(n134), .B(n137), .O(n131));
  invx g100(.A(n133), .O(n132));
  andx g101(.A(n137), .B(n134), .O(n133));
  orx  g102(.A(n135), .B(n170), .O(n134));
  andx g103(.A(n136), .B(pi15), .O(n135));
  andx g104(.A(pi11), .B(n168), .O(n136));
  andx g105(.A(pi14), .B(pi02), .O(n137));
  andx g106(.A(pi13), .B(pi15), .O(n138));
  orx  g107(.A(n140), .B(n177), .O(n139));
  andx g108(.A(n163), .B(n141), .O(n140));
  orx  g109(.A(n142), .B(n181), .O(n141));
  andx g110(.A(pi02), .B(pi12), .O(n142));
  orx  g111(.A(n149), .B(n144), .O(po12));
  andx g112(.A(n146), .B(n145), .O(n144));
  invx g113(.A(n150), .O(n145));
  andx g114(.A(n153), .B(n147), .O(n146));
  invx g115(.A(n148), .O(n147));
  andx g116(.A(n154), .B(n187), .O(n148));
  andx g117(.A(n152), .B(n150), .O(n149));
  orx  g118(.A(n151), .B(n196), .O(n150));
  andx g119(.A(n197), .B(n192), .O(n151));
  invx g120(.A(n153), .O(n152));
  orx  g121(.A(n187), .B(n154), .O(n153));
  andx g122(.A(n156), .B(n155), .O(n154));
  orx  g123(.A(n185), .B(n158), .O(n155));
  invx g124(.A(n157), .O(n156));
  andx g125(.A(n185), .B(n158), .O(n157));
  andx g126(.A(n161), .B(n159), .O(n158));
  invx g127(.A(n160), .O(n159));
  andx g128(.A(n162), .B(n176), .O(n160));
  orx  g129(.A(n176), .B(n162), .O(n161));
  invx g130(.A(n163), .O(n162));
  andx g131(.A(n165), .B(n164), .O(n163));
  orx  g132(.A(n167), .B(n175), .O(n164));
  invx g133(.A(n166), .O(n165));
  andx g134(.A(n175), .B(n167), .O(n166));
  andx g135(.A(n169), .B(n168), .O(n167));
  orx  g136(.A(n171), .B(n174), .O(n168));
  invx g137(.A(n170), .O(n169));
  andx g138(.A(n174), .B(n171), .O(n170));
  orx  g139(.A(n172), .B(n218), .O(n171));
  andx g140(.A(n173), .B(pi15), .O(n172));
  andx g141(.A(pi09), .B(n216), .O(n173));
  andx g142(.A(pi13), .B(pi14), .O(n174));
  andx g143(.A(pi11), .B(pi15), .O(n175));
  orx  g144(.A(n178), .B(n177), .O(n176));
  andx g145(.A(n181), .B(pi02), .O(n177));
  andx g146(.A(n180), .B(n179), .O(n178));
  orx  g147(.A(n720), .B(n303), .O(n179));
  invx g148(.A(n181), .O(n180));
  orx  g149(.A(n182), .B(n225), .O(n181));
  andx g150(.A(n209), .B(n183), .O(n182));
  orx  g151(.A(n184), .B(n229), .O(n183));
  andx g152(.A(pi13), .B(pi12), .O(n184));
  orx  g153(.A(n186), .B(n235), .O(n185));
  andx g154(.A(n206), .B(n232), .O(n186));
  andx g155(.A(n239), .B(n201), .O(n187));
  andx g156(.A(n191), .B(n189), .O(po11));
  invx g157(.A(n190), .O(n189));
  andx g158(.A(n192), .B(n194), .O(n190));
  orx  g159(.A(n194), .B(n192), .O(n191));
  orx  g160(.A(n193), .B(n249), .O(n192));
  andx g161(.A(n312), .B(n251), .O(n193));
  andx g162(.A(n197), .B(n195), .O(n194));
  invx g163(.A(n196), .O(n195));
  andx g164(.A(n198), .B(n255), .O(n196));
  orx  g165(.A(n255), .B(n198), .O(n197));
  orx  g166(.A(n200), .B(n199), .O(n198));
  andx g167(.A(n202), .B(n239), .O(n199));
  andx g168(.A(n238), .B(n201), .O(n200));
  invx g169(.A(n202), .O(n201));
  orx  g170(.A(n205), .B(n203), .O(n202));
  invx g171(.A(n204), .O(n203));
  orx  g172(.A(n206), .B(n231), .O(n204));
  andx g173(.A(n231), .B(n206), .O(n205));
  andx g174(.A(n210), .B(n207), .O(n206));
  orx  g175(.A(n209), .B(n208), .O(n207));
  invx g176(.A(n224), .O(n208));
  invx g177(.A(n211), .O(n209));
  orx  g178(.A(n224), .B(n211), .O(n210));
  orx  g179(.A(n214), .B(n212), .O(n211));
  invx g180(.A(n213), .O(n212));
  orx  g181(.A(n215), .B(n223), .O(n213));
  andx g182(.A(n223), .B(n215), .O(n214));
  andx g183(.A(n217), .B(n216), .O(n215));
  orx  g184(.A(n219), .B(n222), .O(n216));
  invx g185(.A(n218), .O(n217));
  andx g186(.A(n222), .B(n219), .O(n218));
  orx  g187(.A(n220), .B(n276), .O(n219));
  andx g188(.A(n221), .B(pi15), .O(n220));
  andx g189(.A(pi07), .B(n274), .O(n221));
  andx g190(.A(pi11), .B(pi14), .O(n222));
  andx g191(.A(pi09), .B(pi15), .O(n223));
  orx  g192(.A(n226), .B(n225), .O(n224));
  andx g193(.A(n229), .B(pi13), .O(n225));
  andx g194(.A(n228), .B(n227), .O(n226));
  orx  g195(.A(n720), .B(n525), .O(n227));
  invx g196(.A(n229), .O(n228));
  orx  g197(.A(n230), .B(n285), .O(n229));
  andx g198(.A(n269), .B(n286), .O(n230));
  andx g199(.A(n234), .B(n232), .O(n231));
  orx  g200(.A(n233), .B(n236), .O(n232));
  andx g201(.A(pi02), .B(pi10), .O(n233));
  invx g202(.A(n235), .O(n234));
  andx g203(.A(n236), .B(pi02), .O(n235));
  orx  g204(.A(n237), .B(n296), .O(n236));
  andx g205(.A(n265), .B(n293), .O(n237));
  invx g206(.A(n239), .O(n238));
  orx  g207(.A(n240), .B(n300), .O(n239));
  andx g208(.A(n261), .B(n241), .O(n240));
  orx  g209(.A(n242), .B(n305), .O(n241));
  andx g210(.A(pi02), .B(pi08), .O(n242));
  orx  g211(.A(n247), .B(n244), .O(po10));
  andx g212(.A(n246), .B(n245), .O(n244));
  invx g213(.A(n312), .O(n245));
  invx g214(.A(n248), .O(n246));
  andx g215(.A(n312), .B(n248), .O(n247));
  orx  g216(.A(n250), .B(n249), .O(n248));
  andx g217(.A(n252), .B(n311), .O(n249));
  invx g218(.A(n251), .O(n250));
  orx  g219(.A(n311), .B(n252), .O(n251));
  andx g220(.A(n254), .B(n253), .O(n252));
  orx  g221(.A(n309), .B(n256), .O(n253));
  invx g222(.A(n255), .O(n254));
  andx g223(.A(n309), .B(n256), .O(n255));
  andx g224(.A(n259), .B(n257), .O(n256));
  invx g225(.A(n258), .O(n257));
  andx g226(.A(n260), .B(n299), .O(n258));
  orx  g227(.A(n299), .B(n260), .O(n259));
  invx g228(.A(n261), .O(n260));
  andx g229(.A(n263), .B(n262), .O(n261));
  orx  g230(.A(n265), .B(n292), .O(n262));
  invx g231(.A(n264), .O(n263));
  andx g232(.A(n292), .B(n265), .O(n264));
  andx g233(.A(n267), .B(n266), .O(n265));
  orx  g234(.A(n269), .B(n283), .O(n266));
  invx g235(.A(n268), .O(n267));
  andx g236(.A(n283), .B(n269), .O(n268));
  andx g237(.A(n271), .B(n270), .O(n269));
  orx  g238(.A(n273), .B(n282), .O(n270));
  invx g239(.A(n272), .O(n271));
  andx g240(.A(n282), .B(n273), .O(n272));
  andx g241(.A(n275), .B(n274), .O(n273));
  orx  g242(.A(n277), .B(n281), .O(n274));
  invx g243(.A(n276), .O(n275));
  andx g244(.A(n281), .B(n277), .O(n276));
  orx  g245(.A(n279), .B(n278), .O(n277));
  andx g246(.A(n346), .B(n344), .O(n278));
  andx g247(.A(n280), .B(pi14), .O(n279));
  andx g248(.A(pi07), .B(n341), .O(n280));
  andx g249(.A(pi09), .B(pi14), .O(n281));
  andx g250(.A(pi07), .B(pi15), .O(n282));
  andx g251(.A(n286), .B(n284), .O(n283));
  invx g252(.A(n285), .O(n284));
  andx g253(.A(n288), .B(pi11), .O(n285));
  orx  g254(.A(n288), .B(n287), .O(n286));
  andx g255(.A(pi11), .B(pi12), .O(n287));
  orx  g256(.A(n289), .B(n349), .O(n288));
  andx g257(.A(n334), .B(n290), .O(n289));
  orx  g258(.A(n291), .B(n353), .O(n290));
  andx g259(.A(pi12), .B(pi09), .O(n291));
  andx g260(.A(n295), .B(n293), .O(n292));
  orx  g261(.A(n294), .B(n297), .O(n293));
  andx g262(.A(pi13), .B(pi10), .O(n294));
  invx g263(.A(n296), .O(n295));
  andx g264(.A(n297), .B(pi13), .O(n296));
  orx  g265(.A(n298), .B(n359), .O(n297));
  andx g266(.A(n331), .B(n356), .O(n298));
  orx  g267(.A(n301), .B(n300), .O(n299));
  andx g268(.A(n305), .B(pi02), .O(n300));
  andx g269(.A(n304), .B(n302), .O(n301));
  orx  g270(.A(n689), .B(n303), .O(n302));
  invx g271(.A(pi02), .O(n303));
  invx g272(.A(n305), .O(n304));
  orx  g273(.A(n306), .B(n363), .O(n305));
  andx g274(.A(n325), .B(n307), .O(n306));
  orx  g275(.A(n308), .B(n367), .O(n307));
  andx g276(.A(pi13), .B(pi08), .O(n308));
  orx  g277(.A(n310), .B(n373), .O(n309));
  andx g278(.A(n322), .B(n370), .O(n310));
  andx g279(.A(n379), .B(n317), .O(n311));
  andx g280(.A(n460), .B(n313), .O(n312));
  andx g281(.A(n381), .B(n314), .O(n313));
  orx  g282(.A(n316), .B(n315), .O(n314));
  andx g283(.A(n318), .B(n379), .O(n315));
  andx g284(.A(n378), .B(n317), .O(n316));
  invx g285(.A(n318), .O(n317));
  orx  g286(.A(n321), .B(n319), .O(n318));
  invx g287(.A(n320), .O(n319));
  orx  g288(.A(n322), .B(n369), .O(n320));
  andx g289(.A(n369), .B(n322), .O(n321));
  andx g290(.A(n326), .B(n323), .O(n322));
  orx  g291(.A(n325), .B(n324), .O(n323));
  invx g292(.A(n362), .O(n324));
  invx g293(.A(n327), .O(n325));
  orx  g294(.A(n362), .B(n327), .O(n326));
  orx  g295(.A(n330), .B(n328), .O(n327));
  invx g296(.A(n329), .O(n328));
  orx  g297(.A(n331), .B(n355), .O(n329));
  andx g298(.A(n355), .B(n331), .O(n330));
  andx g299(.A(n335), .B(n332), .O(n331));
  orx  g300(.A(n334), .B(n333), .O(n332));
  invx g301(.A(n348), .O(n333));
  invx g302(.A(n336), .O(n334));
  orx  g303(.A(n348), .B(n336), .O(n335));
  orx  g304(.A(n339), .B(n337), .O(n336));
  invx g305(.A(n338), .O(n337));
  orx  g306(.A(n340), .B(n347), .O(n338));
  andx g307(.A(n347), .B(n340), .O(n339));
  andx g308(.A(n342), .B(n341), .O(n340));
  orx  g309(.A(n346), .B(n344), .O(n341));
  orx  g310(.A(n503), .B(n343), .O(n342));
  invx g311(.A(n344), .O(n343));
  orx  g312(.A(n345), .B(n501), .O(n344));
  andx g313(.A(n346), .B(n617), .O(n345));
  invx g314(.A(n503), .O(n346));
  andx g315(.A(pi07), .B(pi14), .O(n347));
  orx  g316(.A(n350), .B(n349), .O(n348));
  andx g317(.A(n353), .B(pi09), .O(n349));
  andx g318(.A(n352), .B(n351), .O(n350));
  orx  g319(.A(n631), .B(n720), .O(n351));
  invx g320(.A(n353), .O(n352));
  orx  g321(.A(n354), .B(n486), .O(n353));
  andx g322(.A(n483), .B(n491), .O(n354));
  andx g323(.A(n358), .B(n356), .O(n355));
  orx  g324(.A(n357), .B(n360), .O(n356));
  andx g325(.A(pi11), .B(pi10), .O(n357));
  invx g326(.A(n359), .O(n358));
  andx g327(.A(n360), .B(pi11), .O(n359));
  orx  g328(.A(n361), .B(n507), .O(n360));
  andx g329(.A(n478), .B(n508), .O(n361));
  orx  g330(.A(n364), .B(n363), .O(n362));
  andx g331(.A(n367), .B(pi13), .O(n363));
  andx g332(.A(n366), .B(n365), .O(n364));
  orx  g333(.A(n689), .B(n525), .O(n365));
  invx g334(.A(n367), .O(n366));
  orx  g335(.A(n368), .B(n516), .O(n367));
  andx g336(.A(n474), .B(n513), .O(n368));
  andx g337(.A(n372), .B(n370), .O(n369));
  orx  g338(.A(n371), .B(n374), .O(n370));
  andx g339(.A(pi02), .B(pi05), .O(n371));
  invx g340(.A(n373), .O(n372));
  andx g341(.A(n374), .B(pi02), .O(n373));
  orx  g342(.A(n375), .B(n522), .O(n374));
  andx g343(.A(n468), .B(n376), .O(n375));
  orx  g344(.A(n377), .B(n527), .O(n376));
  andx g345(.A(pi13), .B(pi05), .O(n377));
  invx g346(.A(n379), .O(n378));
  orx  g347(.A(n380), .B(n533), .O(n379));
  andx g348(.A(n465), .B(n530), .O(n380));
  orx  g349(.A(n383), .B(n382), .O(n381));
  andx g350(.A(n385), .B(pi02), .O(n382));
  andx g351(.A(n451), .B(n384), .O(n383));
  orx  g352(.A(n450), .B(n385), .O(n384));
  orx  g353(.A(n387), .B(n386), .O(n385));
  andx g354(.A(n389), .B(pi13), .O(n386));
  andx g355(.A(n443), .B(n388), .O(n387));
  orx  g356(.A(n442), .B(n389), .O(n388));
  orx  g357(.A(n391), .B(n390), .O(n389));
  andx g358(.A(n393), .B(pi11), .O(n390));
  andx g359(.A(n434), .B(n392), .O(n391));
  orx  g360(.A(n433), .B(n393), .O(n392));
  orx  g361(.A(n395), .B(n394), .O(n393));
  andx g362(.A(n397), .B(pi09), .O(n394));
  andx g363(.A(n427), .B(n396), .O(n395));
  orx  g364(.A(n426), .B(n397), .O(n396));
  invx g365(.A(n398), .O(n397));
  andx g366(.A(n400), .B(n399), .O(n398));
  orx  g367(.A(n402), .B(n416), .O(n399));
  orx  g368(.A(n417), .B(n401), .O(n400));
  andx g369(.A(n414), .B(n402), .O(n401));
  andx g370(.A(n404), .B(n403), .O(n402));
  orx  g371(.A(n410), .B(n406), .O(n403));
  orx  g372(.A(n412), .B(n405), .O(n404));
  andx g373(.A(n410), .B(n406), .O(n405));
  andx g374(.A(n409), .B(n407), .O(n406));
  orx  g375(.A(n408), .B(n661), .O(n407));
  invx g376(.A(n561), .O(n408));
  orx  g377(.A(n660), .B(n561), .O(n409));
  invx g378(.A(n411), .O(n410));
  andx g379(.A(n561), .B(po00), .O(n411));
  invx g380(.A(n413), .O(n412));
  andx g381(.A(pi06), .B(pi01), .O(n413));
  orx  g382(.A(n416), .B(n415), .O(n414));
  invx g383(.A(pi01), .O(n415));
  invx g384(.A(pi07), .O(n416));
  andx g385(.A(n419), .B(n418), .O(n417));
  orx  g386(.A(n421), .B(n554), .O(n418));
  invx g387(.A(n420), .O(n419));
  andx g388(.A(n554), .B(n421), .O(n420));
  andx g389(.A(n423), .B(n422), .O(n421));
  orx  g390(.A(n425), .B(n559), .O(n422));
  invx g391(.A(n424), .O(n423));
  andx g392(.A(n559), .B(n425), .O(n424));
  invx g393(.A(n560), .O(n425));
  andx g394(.A(pi09), .B(pi01), .O(n426));
  orx  g395(.A(n429), .B(n428), .O(n427));
  andx g396(.A(n563), .B(n431), .O(n428));
  invx g397(.A(n430), .O(n429));
  orx  g398(.A(n431), .B(n563), .O(n430));
  orx  g399(.A(n547), .B(n432), .O(n431));
  invx g400(.A(n549), .O(n432));
  andx g401(.A(pi11), .B(pi01), .O(n433));
  orx  g402(.A(n436), .B(n435), .O(n434));
  andx g403(.A(n572), .B(n438), .O(n435));
  invx g404(.A(n437), .O(n436));
  orx  g405(.A(n438), .B(n572), .O(n437));
  orx  g406(.A(n439), .B(n543), .O(n438));
  andx g407(.A(n441), .B(n440), .O(n439));
  orx  g408(.A(n458), .B(n631), .O(n440));
  invx g409(.A(n546), .O(n441));
  andx g410(.A(pi13), .B(pi01), .O(n442));
  invx g411(.A(n444), .O(n443));
  orx  g412(.A(n447), .B(n445), .O(n444));
  invx g413(.A(n446), .O(n445));
  orx  g414(.A(n579), .B(n448), .O(n446));
  andx g415(.A(n448), .B(n579), .O(n447));
  andx g416(.A(n449), .B(n541), .O(n448));
  invx g417(.A(n539), .O(n449));
  andx g418(.A(pi02), .B(pi01), .O(n450));
  orx  g419(.A(n453), .B(n452), .O(n451));
  andx g420(.A(n589), .B(n455), .O(n452));
  invx g421(.A(n454), .O(n453));
  orx  g422(.A(n455), .B(n589), .O(n454));
  orx  g423(.A(n456), .B(n535), .O(n455));
  andx g424(.A(n459), .B(n457), .O(n456));
  orx  g425(.A(n458), .B(n525), .O(n457));
  invx g426(.A(pi03), .O(n458));
  invx g427(.A(n538), .O(n459));
  invx g428(.A(n461), .O(n460));
  orx  g429(.A(n464), .B(n462), .O(n461));
  invx g430(.A(n463), .O(n462));
  orx  g431(.A(n465), .B(n529), .O(n463));
  andx g432(.A(n529), .B(n465), .O(n464));
  andx g433(.A(n469), .B(n466), .O(n465));
  orx  g434(.A(n468), .B(n467), .O(n466));
  invx g435(.A(n521), .O(n467));
  invx g436(.A(n470), .O(n468));
  orx  g437(.A(n521), .B(n470), .O(n469));
  orx  g438(.A(n473), .B(n471), .O(n470));
  invx g439(.A(n472), .O(n471));
  orx  g440(.A(n474), .B(n512), .O(n472));
  andx g441(.A(n512), .B(n474), .O(n473));
  andx g442(.A(n476), .B(n475), .O(n474));
  orx  g443(.A(n478), .B(n505), .O(n475));
  invx g444(.A(n477), .O(n476));
  andx g445(.A(n505), .B(n478), .O(n477));
  andx g446(.A(n481), .B(n479), .O(n478));
  invx g447(.A(n480), .O(n479));
  andx g448(.A(n482), .B(n491), .O(n480));
  orx  g449(.A(n491), .B(n482), .O(n481));
  andx g450(.A(n485), .B(n483), .O(n482));
  orx  g451(.A(n484), .B(n487), .O(n483));
  andx g452(.A(pi12), .B(pi07), .O(n484));
  invx g453(.A(n486), .O(n485));
  andx g454(.A(n487), .B(pi07), .O(n486));
  orx  g455(.A(n489), .B(n488), .O(n487));
  andx g456(.A(n610), .B(n612), .O(n488));
  andx g457(.A(n607), .B(n490), .O(n489));
  orx  g458(.A(n610), .B(n612), .O(n490));
  orx  g459(.A(n494), .B(n492), .O(n491));
  andx g460(.A(n493), .B(n497), .O(n492));
  orx  g461(.A(n721), .B(n504), .O(n493));
  invx g462(.A(n495), .O(n494));
  orx  g463(.A(n496), .B(n721), .O(n495));
  orx  g464(.A(n499), .B(n497), .O(n496));
  andx g465(.A(pi14), .B(n498), .O(n497));
  andx g466(.A(n502), .B(pi06), .O(n498));
  andx g467(.A(n503), .B(n500), .O(n499));
  orx  g468(.A(n504), .B(n501), .O(n500));
  invx g469(.A(n502), .O(n501));
  orx  g470(.A(n614), .B(n616), .O(n502));
  orx  g471(.A(n690), .B(n504), .O(n503));
  invx g472(.A(pi15), .O(n504));
  andx g473(.A(n508), .B(n506), .O(n505));
  invx g474(.A(n507), .O(n506));
  andx g475(.A(n509), .B(pi09), .O(n507));
  orx  g476(.A(n511), .B(n509), .O(n508));
  orx  g477(.A(n510), .B(n623), .O(n509));
  andx g478(.A(n601), .B(n621), .O(n510));
  andx g479(.A(pi10), .B(pi09), .O(n511));
  andx g480(.A(n515), .B(n513), .O(n512));
  orx  g481(.A(n514), .B(n517), .O(n513));
  andx g482(.A(pi11), .B(pi08), .O(n514));
  invx g483(.A(n516), .O(n515));
  andx g484(.A(n517), .B(pi11), .O(n516));
  orx  g485(.A(n518), .B(n628), .O(n517));
  andx g486(.A(n597), .B(n519), .O(n518));
  orx  g487(.A(n520), .B(n633), .O(n519));
  andx g488(.A(pi09), .B(pi08), .O(n520));
  orx  g489(.A(n523), .B(n522), .O(n521));
  andx g490(.A(n527), .B(pi13), .O(n522));
  andx g491(.A(n526), .B(n524), .O(n523));
  orx  g492(.A(n586), .B(n525), .O(n524));
  invx g493(.A(pi13), .O(n525));
  invx g494(.A(n527), .O(n526));
  orx  g495(.A(n528), .B(n639), .O(n527));
  andx g496(.A(n593), .B(n637), .O(n528));
  andx g497(.A(n532), .B(n530), .O(n529));
  orx  g498(.A(n531), .B(n534), .O(n530));
  andx g499(.A(pi02), .B(pi03), .O(n531));
  invx g500(.A(n533), .O(n532));
  andx g501(.A(n534), .B(pi02), .O(n533));
  orx  g502(.A(n536), .B(n535), .O(n534));
  andx g503(.A(n538), .B(pi13), .O(n535));
  andx g504(.A(n589), .B(n537), .O(n536));
  orx  g505(.A(n588), .B(n538), .O(n537));
  orx  g506(.A(n540), .B(n539), .O(n538));
  andx g507(.A(n542), .B(pi11), .O(n539));
  andx g508(.A(n579), .B(n541), .O(n540));
  orx  g509(.A(n578), .B(n542), .O(n541));
  orx  g510(.A(n544), .B(n543), .O(n542));
  andx g511(.A(n546), .B(pi09), .O(n543));
  andx g512(.A(n572), .B(n545), .O(n544));
  orx  g513(.A(n571), .B(n546), .O(n545));
  orx  g514(.A(n548), .B(n547), .O(n546));
  andx g515(.A(n550), .B(pi07), .O(n547));
  andx g516(.A(n563), .B(n549), .O(n548));
  orx  g517(.A(n562), .B(n550), .O(n549));
  orx  g518(.A(n552), .B(n551), .O(n550));
  andx g519(.A(n559), .B(n554), .O(n551));
  andx g520(.A(n560), .B(n553), .O(n552));
  orx  g521(.A(n559), .B(n554), .O(n553));
  orx  g522(.A(n557), .B(n555), .O(n554));
  invx g523(.A(n556), .O(n555));
  orx  g524(.A(n558), .B(n686), .O(n556));
  andx g525(.A(n686), .B(n558), .O(n557));
  orx  g526(.A(n721), .B(n586), .O(n558));
  andx g527(.A(pi06), .B(pi03), .O(n559));
  andx g528(.A(n561), .B(n661), .O(n560));
  andx g529(.A(pi04), .B(pi03), .O(n561));
  andx g530(.A(pi07), .B(pi03), .O(n562));
  orx  g531(.A(n566), .B(n564), .O(n563));
  invx g532(.A(n565), .O(n564));
  orx  g533(.A(n567), .B(n652), .O(n565));
  andx g534(.A(n652), .B(n567), .O(n566));
  andx g535(.A(n570), .B(n568), .O(n567));
  orx  g536(.A(n569), .B(n657), .O(n568));
  invx g537(.A(n656), .O(n569));
  orx  g538(.A(n658), .B(n656), .O(n570));
  andx g539(.A(pi09), .B(pi03), .O(n571));
  orx  g540(.A(n574), .B(n573), .O(n572));
  andx g541(.A(n663), .B(n576), .O(n573));
  invx g542(.A(n575), .O(n574));
  orx  g543(.A(n576), .B(n663), .O(n575));
  orx  g544(.A(n645), .B(n577), .O(n576));
  invx g545(.A(n647), .O(n577));
  andx g546(.A(pi11), .B(pi03), .O(n578));
  andx g547(.A(n582), .B(n580), .O(n579));
  orx  g548(.A(n672), .B(n581), .O(n580));
  invx g549(.A(n583), .O(n581));
  orx  g550(.A(n583), .B(n673), .O(n582));
  orx  g551(.A(n584), .B(n641), .O(n583));
  andx g552(.A(n587), .B(n585), .O(n584));
  orx  g553(.A(n586), .B(n631), .O(n585));
  invx g554(.A(pi05), .O(n586));
  invx g555(.A(n644), .O(n587));
  andx g556(.A(pi13), .B(pi03), .O(n588));
  orx  g557(.A(n591), .B(n590), .O(n589));
  andx g558(.A(n593), .B(n635), .O(n590));
  invx g559(.A(n592), .O(n591));
  orx  g560(.A(n635), .B(n593), .O(n592));
  orx  g561(.A(n595), .B(n594), .O(n593));
  andx g562(.A(n597), .B(n627), .O(n594));
  invx g563(.A(n596), .O(n595));
  orx  g564(.A(n627), .B(n597), .O(n596));
  orx  g565(.A(n599), .B(n598), .O(n597));
  andx g566(.A(n601), .B(n619), .O(n598));
  invx g567(.A(n600), .O(n599));
  orx  g568(.A(n619), .B(n601), .O(n600));
  orx  g569(.A(n604), .B(n602), .O(n601));
  invx g570(.A(n603), .O(n602));
  orx  g571(.A(n605), .B(n612), .O(n603));
  andx g572(.A(n612), .B(n605), .O(n604));
  andx g573(.A(n609), .B(n606), .O(n605));
  orx  g574(.A(n608), .B(n607), .O(n606));
  invx g575(.A(n611), .O(n607));
  invx g576(.A(n610), .O(n608));
  orx  g577(.A(n611), .B(n610), .O(n609));
  andx g578(.A(pi06), .B(pi12), .O(n610));
  orx  g579(.A(n719), .B(n715), .O(n611));
  orx  g580(.A(n615), .B(n613), .O(n612));
  andx g581(.A(n617), .B(n614), .O(n613));
  invx g582(.A(n618), .O(n614));
  andx g583(.A(n618), .B(n616), .O(n615));
  invx g584(.A(n617), .O(n616));
  andx g585(.A(pi04), .B(pi14), .O(n617));
  andx g586(.A(pi00), .B(pi15), .O(n618));
  orx  g587(.A(n623), .B(n620), .O(n619));
  invx g588(.A(n621), .O(n620));
  orx  g589(.A(n622), .B(n624), .O(n621));
  andx g590(.A(pi10), .B(pi07), .O(n622));
  andx g591(.A(n624), .B(pi07), .O(n623));
  orx  g592(.A(n626), .B(n625), .O(n624));
  andx g593(.A(n717), .B(n712), .O(n625));
  andx g594(.A(n723), .B(n711), .O(n626));
  orx  g595(.A(n629), .B(n628), .O(n627));
  andx g596(.A(n633), .B(pi09), .O(n628));
  andx g597(.A(n632), .B(n630), .O(n629));
  orx  g598(.A(n689), .B(n631), .O(n630));
  invx g599(.A(pi09), .O(n631));
  invx g600(.A(n633), .O(n632));
  orx  g601(.A(n634), .B(n679), .O(n633));
  andx g602(.A(n680), .B(n699), .O(n634));
  orx  g603(.A(n639), .B(n636), .O(n635));
  invx g604(.A(n637), .O(n636));
  orx  g605(.A(n638), .B(n640), .O(n637));
  andx g606(.A(pi11), .B(pi05), .O(n638));
  andx g607(.A(n640), .B(pi11), .O(n639));
  orx  g608(.A(n642), .B(n641), .O(n640));
  andx g609(.A(n644), .B(pi09), .O(n641));
  andx g610(.A(n672), .B(n643), .O(n642));
  orx  g611(.A(n671), .B(n644), .O(n643));
  orx  g612(.A(n646), .B(n645), .O(n644));
  andx g613(.A(n648), .B(pi07), .O(n645));
  andx g614(.A(n663), .B(n647), .O(n646));
  orx  g615(.A(n662), .B(n648), .O(n647));
  orx  g616(.A(n650), .B(n649), .O(n648));
  andx g617(.A(n656), .B(n652), .O(n649));
  andx g618(.A(n657), .B(n651), .O(n650));
  orx  g619(.A(n656), .B(n652), .O(n651));
  orx  g620(.A(n655), .B(n653), .O(n652));
  invx g621(.A(n654), .O(n653));
  orx  g622(.A(n659), .B(n722), .O(n654));
  andx g623(.A(n722), .B(n659), .O(n655));
  andx g624(.A(pi06), .B(pi05), .O(n656));
  invx g625(.A(n658), .O(n657));
  orx  g626(.A(n660), .B(n659), .O(n658));
  orx  g627(.A(n721), .B(n689), .O(n659));
  invx g628(.A(n661), .O(n660));
  andx g629(.A(pi00), .B(pi05), .O(n661));
  andx g630(.A(pi07), .B(pi05), .O(n662));
  orx  g631(.A(n666), .B(n664), .O(n663));
  invx g632(.A(n665), .O(n664));
  orx  g633(.A(n667), .B(n691), .O(n665));
  andx g634(.A(n691), .B(n667), .O(n666));
  andx g635(.A(n669), .B(n668), .O(n667));
  orx  g636(.A(n688), .B(n685), .O(n668));
  invx g637(.A(n670), .O(n669));
  andx g638(.A(n685), .B(n688), .O(n670));
  andx g639(.A(pi09), .B(pi05), .O(n671));
  invx g640(.A(n673), .O(n672));
  orx  g641(.A(n675), .B(n674), .O(n673));
  andx g642(.A(n677), .B(n699), .O(n674));
  invx g643(.A(n676), .O(n675));
  orx  g644(.A(n699), .B(n677), .O(n676));
  andx g645(.A(n680), .B(n678), .O(n677));
  invx g646(.A(n679), .O(n678));
  andx g647(.A(n681), .B(pi07), .O(n679));
  orx  g648(.A(n698), .B(n681), .O(n680));
  orx  g649(.A(n683), .B(n682), .O(n681));
  andx g650(.A(n687), .B(n685), .O(n682));
  andx g651(.A(n691), .B(n684), .O(n683));
  orx  g652(.A(n687), .B(n685), .O(n684));
  andx g653(.A(n686), .B(n697), .O(n685));
  andx g654(.A(pi00), .B(pi08), .O(n686));
  invx g655(.A(n688), .O(n687));
  orx  g656(.A(n690), .B(n689), .O(n688));
  invx g657(.A(pi08), .O(n689));
  invx g658(.A(pi06), .O(n690));
  orx  g659(.A(n693), .B(n692), .O(n691));
  andx g660(.A(n695), .B(n696), .O(n692));
  invx g661(.A(n694), .O(n693));
  orx  g662(.A(n696), .B(n695), .O(n694));
  andx g663(.A(pi00), .B(pi12), .O(n695));
  invx g664(.A(n697), .O(n696));
  andx g665(.A(pi04), .B(pi10), .O(n697));
  andx g666(.A(pi08), .B(pi07), .O(n698));
  orx  g667(.A(n709), .B(n700), .O(n699));
  orx  g668(.A(n703), .B(n701), .O(n700));
  invx g669(.A(n702), .O(n701));
  orx  g670(.A(n704), .B(n712), .O(n702));
  andx g671(.A(n705), .B(n704), .O(n703));
  orx  g672(.A(n723), .B(n708), .O(n704));
  andx g673(.A(n712), .B(n706), .O(n705));
  invx g674(.A(n707), .O(n706));
  andx g675(.A(n708), .B(n723), .O(n707));
  invx g676(.A(n717), .O(n708));
  andx g677(.A(n723), .B(n710), .O(n709));
  invx g678(.A(n711), .O(n710));
  orx  g679(.A(n717), .B(n712), .O(n711));
  orx  g680(.A(n714), .B(n713), .O(n712));
  andx g681(.A(n716), .B(n719), .O(n713));
  andx g682(.A(n718), .B(n715), .O(n714));
  invx g683(.A(n716), .O(n715));
  andx g684(.A(pi00), .B(pi14), .O(n716));
  andx g685(.A(n722), .B(n718), .O(n717));
  invx g686(.A(n719), .O(n718));
  orx  g687(.A(n721), .B(n720), .O(n719));
  invx g688(.A(pi12), .O(n720));
  invx g689(.A(pi04), .O(n721));
  andx g690(.A(pi00), .B(pi10), .O(n722));
  andx g691(.A(pi06), .B(pi10), .O(n723));
  andx g692(.A(pi01), .B(pi00), .O(po00));
endmodule


