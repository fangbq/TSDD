// Benchmark "cosin" written by ABC on Fri Feb  7 13:42:00 2014

module cosin ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63;
  wire n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
    n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
    n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
    n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
    n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
    n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750;
  bufx g0000(.A(n2725), .O(po00));
  bufx g0001(.A(n2724), .O(po01));
  bufx g0002(.A(n2723), .O(po02));
  bufx g0003(.A(n2722), .O(po03));
  bufx g0004(.A(n2721), .O(po04));
  bufx g0005(.A(n2720), .O(po05));
  bufx g0006(.A(n2719), .O(po06));
  bufx g0007(.A(n2718), .O(po07));
  bufx g0008(.A(n2717), .O(po08));
  bufx g0009(.A(n2716), .O(po09));
  bufx g0010(.A(n2715), .O(po10));
  bufx g0011(.A(n2714), .O(po11));
  bufx g0012(.A(n2713), .O(po12));
  bufx g0013(.A(n2712), .O(po13));
  bufx g0014(.A(n2711), .O(po14));
  bufx g0015(.A(n2710), .O(po15));
  bufx g0016(.A(n2709), .O(po16));
  bufx g0017(.A(n2708), .O(po17));
  bufx g0018(.A(n2707), .O(po18));
  bufx g0019(.A(n2706), .O(po19));
  bufx g0020(.A(n2705), .O(po20));
  bufx g0021(.A(n2704), .O(po21));
  bufx g0022(.A(n2703), .O(po22));
  bufx g0023(.A(n2702), .O(po23));
  bufx g0024(.A(n2701), .O(po24));
  bufx g0025(.A(n2700), .O(po25));
  bufx g0026(.A(n2699), .O(po26));
  bufx g0027(.A(n2698), .O(po27));
  bufx g0028(.A(n2697), .O(po28));
  bufx g0029(.A(n2696), .O(po29));
  bufx g0030(.A(n2695), .O(po30));
  bufx g0031(.A(n2694), .O(po31));
  bufx g0032(.A(n2693), .O(po32));
  bufx g0033(.A(n2692), .O(po33));
  bufx g0034(.A(n2691), .O(po34));
  bufx g0035(.A(n2690), .O(po35));
  bufx g0036(.A(n2689), .O(po36));
  bufx g0037(.A(n2688), .O(po37));
  bufx g0038(.A(n2687), .O(po38));
  bufx g0039(.A(n2686), .O(po39));
  bufx g0040(.A(n2685), .O(po40));
  bufx g0041(.A(n2684), .O(po41));
  bufx g0042(.A(n2683), .O(po42));
  bufx g0043(.A(n2682), .O(po43));
  bufx g0044(.A(n2681), .O(po44));
  bufx g0045(.A(n2680), .O(po45));
  bufx g0046(.A(n2679), .O(po46));
  bufx g0047(.A(n2678), .O(po47));
  bufx g0048(.A(n2677), .O(po48));
  bufx g0049(.A(n2676), .O(po49));
  bufx g0050(.A(n2675), .O(po50));
  bufx g0051(.A(n2674), .O(po51));
  bufx g0052(.A(n2642), .O(po52));
  bufx g0053(.A(n2641), .O(po53));
  bufx g0054(.A(n2640), .O(po54));
  bufx g0055(.A(n2639), .O(po55));
  bufx g0056(.A(n2639), .O(po56));
  bufx g0057(.A(n2639), .O(po57));
  bufx g0058(.A(n2639), .O(po58));
  bufx g0059(.A(n2639), .O(po59));
  bufx g0060(.A(n2639), .O(po60));
  bufx g0061(.A(n2639), .O(po61));
  bufx g0062(.A(n2639), .O(po62));
  bufx g0063(.A(n2625), .O(po63));
  orx  g0064(.A(n2671), .B(pi31), .O(n163));
  orx  g0065(.A(pi29), .B(n2320), .O(n164));
  andx g0066(.A(pi27), .B(n215), .O(n165));
  orx  g0067(.A(pi29), .B(pi31), .O(n166));
  orx  g0068(.A(n2316), .B(pi30), .O(n167));
  andx g0069(.A(n230), .B(pi27), .O(n168));
  orx  g0070(.A(n2559), .B(n2277), .O(n169));
  orx  g0071(.A(n2371), .B(n2291), .O(n170));
  orx  g0072(.A(n2539), .B(n2283), .O(n171));
  andx g0073(.A(n1165), .B(pi28), .O(n172));
  orx  g0074(.A(n2543), .B(n2316), .O(n173));
  andx g0075(.A(n1024), .B(pi27), .O(n174));
  andx g0076(.A(n1165), .B(pi27), .O(n175));
  orx  g0077(.A(n2313), .B(n2409), .O(n176));
  orx  g0078(.A(n2282), .B(pi30), .O(n177));
  andx g0079(.A(n340), .B(n192), .O(n178));
  andx g0080(.A(n617), .B(n2482), .O(n179));
  orx  g0081(.A(n2613), .B(n2303), .O(n180));
  orx  g0082(.A(pi28), .B(n2358), .O(n181));
  andx g0083(.A(n2593), .B(n2464), .O(n182));
  andx g0084(.A(n289), .B(n2464), .O(n183));
  andx g0085(.A(pi25), .B(n879), .O(n184));
  andx g0086(.A(n1025), .B(pi27), .O(n185));
  andx g0087(.A(pi27), .B(n2570), .O(n186));
  andx g0088(.A(pi27), .B(n204), .O(n187));
  andx g0089(.A(n2544), .B(pi26), .O(n188));
  andx g0090(.A(n2527), .B(n2285), .O(n189));
  orx  g0091(.A(n2292), .B(n2319), .O(n190));
  orx  g0092(.A(n2559), .B(n2313), .O(n191));
  orx  g0093(.A(n2318), .B(n2409), .O(n192));
  orx  g0094(.A(n1972), .B(n2409), .O(n193));
  orx  g0095(.A(pi31), .B(pi30), .O(n194));
  orx  g0096(.A(pi30), .B(n2302), .O(n195));
  orx  g0097(.A(pi30), .B(n2314), .O(n196));
  orx  g0098(.A(n2273), .B(n2586), .O(n197));
  orx  g0099(.A(pi30), .B(n2318), .O(n198));
  orx  g0100(.A(pi30), .B(n2317), .O(n199));
  orx  g0101(.A(n2290), .B(n2539), .O(n200));
  orx  g0102(.A(n2282), .B(n2586), .O(n201));
  orx  g0103(.A(pi30), .B(n2290), .O(n202));
  orx  g0104(.A(n2282), .B(n2537), .O(n203));
  orx  g0105(.A(n2276), .B(n2543), .O(n204));
  orx  g0106(.A(n348), .B(n349), .O(n205));
  orx  g0107(.A(n429), .B(n430), .O(n206));
  orx  g0108(.A(n484), .B(n485), .O(n207));
  orx  g0109(.A(n802), .B(n803), .O(n208));
  orx  g0110(.A(n723), .B(n370), .O(n209));
  orx  g0111(.A(n371), .B(n372), .O(n210));
  orx  g0112(.A(n367), .B(n368), .O(n211));
  orx  g0113(.A(n625), .B(n366), .O(n212));
  orx  g0114(.A(n358), .B(n359), .O(n213));
  orx  g0115(.A(n472), .B(n347), .O(n214));
  orx  g0116(.A(n345), .B(n346), .O(n215));
  andx g0117(.A(n373), .B(n2464), .O(n216));
  orx  g0118(.A(n375), .B(n374), .O(n217));
  orx  g0119(.A(n393), .B(n394), .O(n218));
  orx  g0120(.A(n391), .B(n392), .O(n219));
  orx  g0121(.A(n723), .B(n378), .O(n220));
  orx  g0122(.A(n376), .B(n377), .O(n221));
  andx g0123(.A(n397), .B(n2465), .O(n222));
  orx  g0124(.A(n399), .B(n398), .O(n223));
  andx g0125(.A(n400), .B(n1023), .O(n224));
  andx g0126(.A(n418), .B(n2295), .O(n225));
  orx  g0127(.A(n419), .B(n420), .O(n226));
  orx  g0128(.A(n439), .B(n440), .O(n227));
  orx  g0129(.A(n437), .B(n438), .O(n228));
  orx  g0130(.A(n425), .B(n426), .O(n229));
  orx  g0131(.A(n2559), .B(n2303), .O(n230));
  andx g0132(.A(n443), .B(n2465), .O(n231));
  orx  g0133(.A(n445), .B(n444), .O(n232));
  orx  g0134(.A(n472), .B(n473), .O(n233));
  orx  g0135(.A(n469), .B(n470), .O(n234));
  orx  g0136(.A(n467), .B(n468), .O(n235));
  orx  g0137(.A(n447), .B(n448), .O(n236));
  orx  g0138(.A(n457), .B(n458), .O(n237));
  orx  g0139(.A(n451), .B(n452), .O(n238));
  orx  g0140(.A(n1862), .B(n446), .O(n239));
  andx g0141(.A(n475), .B(n2465), .O(n240));
  orx  g0142(.A(n477), .B(n476), .O(n241));
  orx  g0143(.A(n492), .B(n493), .O(n242));
  orx  g0144(.A(n480), .B(n481), .O(n243));
  andx g0145(.A(n501), .B(n2465), .O(n244));
  orx  g0146(.A(n503), .B(n502), .O(n245));
  orx  g0147(.A(n518), .B(n519), .O(n246));
  orx  g0148(.A(n509), .B(n510), .O(n247));
  andx g0149(.A(n521), .B(n2479), .O(n248));
  orx  g0150(.A(n523), .B(n522), .O(n249));
  orx  g0151(.A(n540), .B(n541), .O(n250));
  orx  g0152(.A(n532), .B(n533), .O(n251));
  andx g0153(.A(n2542), .B(n906), .O(n252));
  orx  g0154(.A(n524), .B(n525), .O(n253));
  andx g0155(.A(n543), .B(n2478), .O(n254));
  orx  g0156(.A(n545), .B(n544), .O(n255));
  andx g0157(.A(n336), .B(n1017), .O(n256));
  orx  g0158(.A(n798), .B(n554), .O(n257));
  andx g0159(.A(n1028), .B(n1027), .O(n258));
  andx g0160(.A(n562), .B(n2477), .O(n259));
  orx  g0161(.A(n564), .B(n563), .O(n260));
  orx  g0162(.A(n573), .B(n574), .O(n261));
  andx g0163(.A(n584), .B(n2464), .O(n262));
  orx  g0164(.A(n586), .B(n585), .O(n263));
  orx  g0165(.A(n594), .B(n595), .O(n264));
  orx  g0166(.A(n625), .B(n591), .O(n265));
  andx g0167(.A(n602), .B(n2466), .O(n266));
  orx  g0168(.A(n604), .B(n603), .O(n267));
  andx g0169(.A(n618), .B(n2466), .O(n268));
  andx g0170(.A(n1031), .B(n1030), .O(n269));
  orx  g0171(.A(n622), .B(n621), .O(n270));
  andx g0172(.A(n641), .B(n2466), .O(n271));
  orx  g0173(.A(n643), .B(n642), .O(n272));
  andx g0174(.A(pi30), .B(n2319), .O(n273));
  orx  g0175(.A(n646), .B(n647), .O(n274));
  andx g0176(.A(n662), .B(n2466), .O(n275));
  orx  g0177(.A(n664), .B(n663), .O(n276));
  orx  g0178(.A(n670), .B(n671), .O(n277));
  andx g0179(.A(n682), .B(n2467), .O(n278));
  orx  g0180(.A(n684), .B(n683), .O(n279));
  orx  g0181(.A(n685), .B(n686), .O(n280));
  andx g0182(.A(n706), .B(n2467), .O(n281));
  orx  g0183(.A(n708), .B(n707), .O(n282));
  orx  g0184(.A(n723), .B(n724), .O(n283));
  orx  g0185(.A(n711), .B(n712), .O(n284));
  andx g0186(.A(n341), .B(n1034), .O(n285));
  orx  g0187(.A(n728), .B(n727), .O(n286));
  andx g0188(.A(n2308), .B(n176), .O(n287));
  orx  g0189(.A(n472), .B(n740), .O(n288));
  orx  g0190(.A(n735), .B(n736), .O(n289));
  andx g0191(.A(n1035), .B(n1031), .O(n290));
  andx g0192(.A(n737), .B(n734), .O(n291));
  andx g0193(.A(n743), .B(n2467), .O(n292));
  orx  g0194(.A(n745), .B(n744), .O(n293));
  andx g0195(.A(n342), .B(n763), .O(n294));
  orx  g0196(.A(n765), .B(n764), .O(n295));
  orx  g0197(.A(n774), .B(n775), .O(n296));
  orx  g0198(.A(n768), .B(n769), .O(n297));
  andx g0199(.A(n788), .B(n2467), .O(n298));
  orx  g0200(.A(n790), .B(n789), .O(n299));
  andx g0201(.A(n237), .B(n2468), .O(n300));
  orx  g0202(.A(n798), .B(n799), .O(n301));
  andx g0203(.A(n812), .B(n810), .O(n302));
  orx  g0204(.A(n814), .B(n813), .O(n303));
  andx g0205(.A(n834), .B(n2468), .O(n304));
  orx  g0206(.A(n836), .B(n835), .O(n305));
  orx  g0207(.A(n837), .B(n838), .O(n306));
  andx g0208(.A(n839), .B(n1038), .O(n307));
  andx g0209(.A(n851), .B(n2468), .O(n308));
  orx  g0210(.A(n853), .B(n852), .O(n309));
  andx g0211(.A(n868), .B(n2468), .O(n310));
  orx  g0212(.A(n870), .B(n869), .O(n311));
  andx g0213(.A(n209), .B(n1027), .O(n312));
  orx  g0214(.A(n877), .B(n878), .O(n313));
  andx g0215(.A(n886), .B(n2469), .O(n314));
  orx  g0216(.A(n888), .B(n887), .O(n315));
  andx g0217(.A(n2589), .B(n1018), .O(n316));
  orx  g0218(.A(n898), .B(n899), .O(n317));
  orx  g0219(.A(n889), .B(n890), .O(n318));
  andx g0220(.A(n1041), .B(n193), .O(n319));
  andx g0221(.A(n907), .B(n2469), .O(n320));
  orx  g0222(.A(n909), .B(n908), .O(n321));
  andx g0223(.A(n926), .B(n2469), .O(n322));
  orx  g0224(.A(n928), .B(n927), .O(n323));
  andx g0225(.A(n941), .B(n2469), .O(n324));
  orx  g0226(.A(n943), .B(n942), .O(n325));
  andx g0227(.A(n2529), .B(n1018), .O(n326));
  andx g0228(.A(n959), .B(n2470), .O(n327));
  orx  g0229(.A(n961), .B(n960), .O(n328));
  andx g0230(.A(n2561), .B(n1045), .O(n329));
  andx g0231(.A(n977), .B(n2470), .O(n330));
  orx  g0232(.A(n979), .B(n978), .O(n331));
  andx g0233(.A(n994), .B(n2261), .O(n332));
  orx  g0234(.A(n995), .B(n996), .O(n333));
  andx g0235(.A(n344), .B(n1012), .O(n334));
  orx  g0236(.A(n1013), .B(n1014), .O(n335));
  orx  g0237(.A(n2302), .B(n2408), .O(n336));
  orx  g0238(.A(n2308), .B(n2586), .O(n337));
  orx  g0239(.A(pi30), .B(n2307), .O(n338));
  orx  g0240(.A(pi29), .B(n2408), .O(n339));
  andx g0241(.A(pi27), .B(n2470), .O(n340));
  andx g0242(.A(n726), .B(n2470), .O(n341));
  andx g0243(.A(n1036), .B(n2471), .O(n342));
  orx  g0244(.A(n2428), .B(n2673), .O(n343));
  andx g0245(.A(n1020), .B(n2294), .O(n344));
  andx g0246(.A(n2281), .B(n2379), .O(n345));
  andx g0247(.A(pi30), .B(n2314), .O(n346));
  andx g0248(.A(n2273), .B(n2377), .O(n347));
  andx g0249(.A(pi31), .B(n2671), .O(n348));
  andx g0250(.A(pi29), .B(n2321), .O(n349));
  andx g0251(.A(n2280), .B(n2377), .O(n350));
  andx g0252(.A(n2289), .B(pi30), .O(n351));
  andx g0253(.A(n214), .B(n2339), .O(n352));
  andx g0254(.A(n1047), .B(pi27), .O(n353));
  andx g0255(.A(n1021), .B(n2435), .O(n354));
  andx g0256(.A(n1048), .B(pi28), .O(n355));
  andx g0257(.A(n2583), .B(pi27), .O(n356));
  andx g0258(.A(n167), .B(n2335), .O(n357));
  andx g0259(.A(pi30), .B(pi31), .O(n358));
  andx g0260(.A(n2307), .B(n2378), .O(n359));
  andx g0261(.A(n2560), .B(n2335), .O(n360));
  andx g0262(.A(n213), .B(pi27), .O(n361));
  andx g0263(.A(n1050), .B(n2431), .O(n362));
  andx g0264(.A(n1051), .B(pi28), .O(n363));
  andx g0265(.A(n1049), .B(n2471), .O(n364));
  andx g0266(.A(n1052), .B(pi25), .O(n365));
  andx g0267(.A(pi30), .B(n2283), .O(n366));
  andx g0268(.A(pi29), .B(n2388), .O(n367));
  andx g0269(.A(n2308), .B(pi30), .O(n368));
  andx g0270(.A(n1055), .B(n1054), .O(n369));
  andx g0271(.A(n205), .B(n2377), .O(n370));
  andx g0272(.A(n209), .B(n2335), .O(n371));
  andx g0273(.A(n2523), .B(pi27), .O(n372));
  andx g0274(.A(n1057), .B(n1056), .O(n373));
  andx g0275(.A(n1053), .B(n2287), .O(n374));
  andx g0276(.A(n216), .B(pi26), .O(n375));
  andx g0277(.A(n2307), .B(pi30), .O(n376));
  andx g0278(.A(n166), .B(n2379), .O(n377));
  andx g0279(.A(n2314), .B(n2378), .O(n378));
  andx g0280(.A(n221), .B(n2339), .O(n379));
  andx g0281(.A(n220), .B(pi27), .O(n380));
  andx g0282(.A(n215), .B(pi27), .O(n381));
  andx g0283(.A(n2603), .B(n2335), .O(n382));
  andx g0284(.A(n1058), .B(n2438), .O(n383));
  andx g0285(.A(n1059), .B(pi28), .O(n384));
  andx g0286(.A(n2582), .B(pi27), .O(n385));
  andx g0287(.A(n169), .B(n2336), .O(n386));
  andx g0288(.A(n1022), .B(n2432), .O(n387));
  andx g0289(.A(n1061), .B(pi28), .O(n388));
  andx g0290(.A(n1060), .B(n2471), .O(n389));
  andx g0291(.A(n1062), .B(pi25), .O(n390));
  andx g0292(.A(pi30), .B(pi29), .O(n391));
  andx g0293(.A(pi31), .B(n2378), .O(n392));
  andx g0294(.A(pi30), .B(pi29), .O(n393));
  andx g0295(.A(n2290), .B(n2378), .O(n394));
  andx g0296(.A(n1065), .B(n1064), .O(n395));
  andx g0297(.A(n1067), .B(n1066), .O(n396));
  andx g0298(.A(n1069), .B(n1068), .O(n397));
  andx g0299(.A(n1063), .B(n2260), .O(n398));
  andx g0300(.A(n222), .B(pi26), .O(n399));
  andx g0301(.A(n1071), .B(n1070), .O(n400));
  andx g0302(.A(pi30), .B(n2315), .O(n401));
  andx g0303(.A(n2274), .B(n2379), .O(n402));
  andx g0304(.A(n1072), .B(n2294), .O(n403));
  andx g0305(.A(n2529), .B(pi26), .O(n404));
  andx g0306(.A(n224), .B(n2341), .O(n405));
  andx g0307(.A(n1073), .B(pi27), .O(n406));
  andx g0308(.A(pi26), .B(n2291), .O(n407));
  andx g0309(.A(n2581), .B(n2259), .O(n408));
  andx g0310(.A(n213), .B(n2286), .O(n409));
  andx g0311(.A(n2528), .B(pi26), .O(n410));
  andx g0312(.A(n1075), .B(n2336), .O(n411));
  andx g0313(.A(n1076), .B(pi27), .O(n412));
  andx g0314(.A(n1074), .B(n2435), .O(n413));
  andx g0315(.A(n1077), .B(pi28), .O(n414));
  andx g0316(.A(n1080), .B(n1079), .O(n415));
  andx g0317(.A(n1082), .B(n1081), .O(n416));
  andx g0318(.A(n1084), .B(n1083), .O(n417));
  andx g0319(.A(n1086), .B(n1085), .O(n418));
  andx g0320(.A(n1078), .B(n2471), .O(n419));
  andx g0321(.A(n225), .B(pi25), .O(n420));
  andx g0322(.A(n230), .B(n2336), .O(n421));
  andx g0323(.A(n2527), .B(pi27), .O(n422));
  andx g0324(.A(n1087), .B(n2432), .O(n423));
  andx g0325(.A(pi28), .B(n1016), .O(n424));
  andx g0326(.A(pi30), .B(n164), .O(n425));
  andx g0327(.A(n2289), .B(n2380), .O(n426));
  andx g0328(.A(n2273), .B(pi27), .O(n427));
  andx g0329(.A(n229), .B(n2336), .O(n428));
  andx g0330(.A(pi31), .B(n2380), .O(n429));
  andx g0331(.A(pi30), .B(n2321), .O(n430));
  andx g0332(.A(pi27), .B(n192), .O(n431));
  andx g0333(.A(n2579), .B(n2339), .O(n432));
  andx g0334(.A(n1089), .B(n2438), .O(n433));
  andx g0335(.A(n1090), .B(pi28), .O(n434));
  andx g0336(.A(n1088), .B(n2472), .O(n435));
  andx g0337(.A(n1091), .B(pi25), .O(n436));
  andx g0338(.A(n2308), .B(n2379), .O(n437));
  andx g0339(.A(n2317), .B(pi30), .O(n438));
  andx g0340(.A(pi31), .B(n2380), .O(n439));
  andx g0341(.A(pi30), .B(n2312), .O(n440));
  andx g0342(.A(n1094), .B(n1093), .O(n441));
  andx g0343(.A(n1096), .B(n1095), .O(n442));
  andx g0344(.A(n1098), .B(n1097), .O(n443));
  andx g0345(.A(n1092), .B(n2260), .O(n444));
  andx g0346(.A(n231), .B(pi26), .O(n445));
  andx g0347(.A(n2283), .B(n2380), .O(n446));
  andx g0348(.A(n2669), .B(n2320), .O(n447));
  andx g0349(.A(n2276), .B(pi30), .O(n448));
  andx g0350(.A(n239), .B(n2472), .O(n449));
  andx g0351(.A(n2576), .B(pi25), .O(n450));
  andx g0352(.A(n2303), .B(n2380), .O(n451));
  andx g0353(.A(n2307), .B(pi30), .O(n452));
  andx g0354(.A(pi25), .B(n2283), .O(n453));
  andx g0355(.A(n238), .B(n2472), .O(n454));
  andx g0356(.A(n1099), .B(n2337), .O(n455));
  andx g0357(.A(n1100), .B(pi27), .O(n456));
  andx g0358(.A(n2283), .B(n2381), .O(n457));
  andx g0359(.A(pi30), .B(n2316), .O(n458));
  andx g0360(.A(n237), .B(n2472), .O(n459));
  andx g0361(.A(n170), .B(pi25), .O(n460));
  andx g0362(.A(n236), .B(n2473), .O(n461));
  andx g0363(.A(n1024), .B(pi25), .O(n462));
  andx g0364(.A(n1102), .B(n2337), .O(n463));
  andx g0365(.A(n1103), .B(pi27), .O(n464));
  andx g0366(.A(n1101), .B(n2432), .O(n465));
  andx g0367(.A(n1104), .B(pi28), .O(n466));
  andx g0368(.A(pi31), .B(n2381), .O(n467));
  andx g0369(.A(pi30), .B(n2314), .O(n468));
  andx g0370(.A(n2315), .B(n2381), .O(n469));
  andx g0371(.A(n2317), .B(pi30), .O(n470));
  andx g0372(.A(n1107), .B(n1106), .O(n471));
  andx g0373(.A(pi30), .B(n2291), .O(n472));
  andx g0374(.A(pi31), .B(n2382), .O(n473));
  andx g0375(.A(n1109), .B(n1108), .O(n474));
  andx g0376(.A(n1111), .B(n1110), .O(n475));
  andx g0377(.A(n1105), .B(n2295), .O(n476));
  andx g0378(.A(n240), .B(pi26), .O(n477));
  andx g0379(.A(pi29), .B(n2381), .O(n478));
  andx g0380(.A(pi30), .B(n2313), .O(n479));
  andx g0381(.A(pi30), .B(n2282), .O(n480));
  andx g0382(.A(n2313), .B(n2399), .O(n481));
  andx g0383(.A(n1112), .B(n2337), .O(n482));
  andx g0384(.A(n243), .B(pi27), .O(n483));
  andx g0385(.A(n2308), .B(pi30), .O(n484));
  andx g0386(.A(n205), .B(n2382), .O(n485));
  andx g0387(.A(n2302), .B(n2337), .O(n486));
  andx g0388(.A(n2571), .B(pi27), .O(n487));
  andx g0389(.A(n1113), .B(n2439), .O(n488));
  andx g0390(.A(n1114), .B(pi28), .O(n489));
  andx g0391(.A(n171), .B(n2338), .O(n490));
  andx g0392(.A(n2541), .B(pi27), .O(n491));
  andx g0393(.A(pi29), .B(n2390), .O(n492));
  andx g0394(.A(n2277), .B(pi30), .O(n493));
  andx g0395(.A(n206), .B(pi27), .O(n494));
  andx g0396(.A(n242), .B(n2338), .O(n495));
  andx g0397(.A(n1116), .B(n2432), .O(n496));
  andx g0398(.A(n1117), .B(pi28), .O(n497));
  andx g0399(.A(n1115), .B(n2473), .O(n498));
  andx g0400(.A(n1118), .B(pi25), .O(n499));
  andx g0401(.A(n1121), .B(n1120), .O(n500));
  andx g0402(.A(n1123), .B(n1122), .O(n501));
  andx g0403(.A(n1119), .B(n2633), .O(n502));
  andx g0404(.A(n244), .B(pi26), .O(n503));
  andx g0405(.A(n2603), .B(pi28), .O(n504));
  andx g0406(.A(n239), .B(n2437), .O(n505));
  andx g0407(.A(n1124), .B(n2338), .O(n506));
  andx g0408(.A(n1026), .B(pi27), .O(n507));
  andx g0409(.A(n2277), .B(pi30), .O(n508));
  andx g0410(.A(pi29), .B(n2387), .O(n509));
  andx g0411(.A(pi30), .B(n2282), .O(n510));
  andx g0412(.A(n2578), .B(n2433), .O(n511));
  andx g0413(.A(n247), .B(pi28), .O(n512));
  andx g0414(.A(n1126), .B(n2340), .O(n513));
  andx g0415(.A(n1127), .B(pi27), .O(n514));
  andx g0416(.A(n1125), .B(n2473), .O(n515));
  andx g0417(.A(n1128), .B(pi25), .O(n516));
  andx g0418(.A(n1131), .B(n1130), .O(n517));
  andx g0419(.A(pi30), .B(pi29), .O(n518));
  andx g0420(.A(n2315), .B(n2382), .O(n519));
  andx g0421(.A(n1133), .B(n1132), .O(n520));
  andx g0422(.A(n1135), .B(n1134), .O(n521));
  andx g0423(.A(n1129), .B(n2285), .O(n522));
  andx g0424(.A(n248), .B(pi26), .O(n523));
  andx g0425(.A(pi29), .B(n2384), .O(n524));
  andx g0426(.A(pi30), .B(n2303), .O(n525));
  andx g0427(.A(n2560), .B(n2338), .O(n526));
  andx g0428(.A(n253), .B(pi27), .O(n527));
  andx g0429(.A(n2568), .B(pi27), .O(n528));
  andx g0430(.A(n173), .B(n2340), .O(n529));
  andx g0431(.A(n1136), .B(n2668), .O(n530));
  andx g0432(.A(n1137), .B(pi28), .O(n531));
  andx g0433(.A(n2277), .B(pi30), .O(n532));
  andx g0434(.A(n2290), .B(n2382), .O(n533));
  andx g0435(.A(n2580), .B(pi27), .O(n534));
  andx g0436(.A(n251), .B(n2339), .O(n535));
  andx g0437(.A(n1139), .B(n2433), .O(n536));
  andx g0438(.A(n252), .B(pi28), .O(n537));
  andx g0439(.A(n1138), .B(n2473), .O(n538));
  andx g0440(.A(n1140), .B(pi25), .O(n539));
  andx g0441(.A(n2528), .B(pi27), .O(n540));
  andx g0442(.A(n2525), .B(n2340), .O(n541));
  orx  g0443(.A(n174), .B(n2573), .O(n542));
  andx g0444(.A(n1143), .B(n1142), .O(n543));
  andx g0445(.A(n1141), .B(n2262), .O(n544));
  andx g0446(.A(n254), .B(pi26), .O(n545));
  orx  g0447(.A(n2312), .B(n2539), .O(n546));
  andx g0448(.A(n236), .B(pi27), .O(n547));
  andx g0449(.A(n2540), .B(n2341), .O(n548));
  andx g0450(.A(n1144), .B(n2435), .O(n549));
  andx g0451(.A(n258), .B(pi28), .O(n550));
  andx g0452(.A(n1147), .B(n1146), .O(n551));
  andx g0453(.A(pi27), .B(n2545), .O(n552));
  andx g0454(.A(n551), .B(n2340), .O(n553));
  andx g0455(.A(n2275), .B(n2383), .O(n554));
  andx g0456(.A(n214), .B(pi27), .O(n555));
  andx g0457(.A(n257), .B(n2341), .O(n556));
  andx g0458(.A(n1148), .B(n2433), .O(n557));
  andx g0459(.A(n1149), .B(pi28), .O(n558));
  andx g0460(.A(n1145), .B(n2474), .O(n559));
  andx g0461(.A(n1150), .B(pi25), .O(n560));
  andx g0462(.A(n1153), .B(n1152), .O(n561));
  andx g0463(.A(n1155), .B(n1154), .O(n562));
  andx g0464(.A(n1151), .B(n2294), .O(n563));
  andx g0465(.A(n259), .B(pi26), .O(n564));
  andx g0466(.A(n166), .B(pi27), .O(n565));
  andx g0467(.A(n1158), .B(n1157), .O(n566));
  andx g0468(.A(n1156), .B(n2436), .O(n567));
  andx g0469(.A(n566), .B(pi28), .O(n568));
  andx g0470(.A(pi31), .B(n2383), .O(n569));
  andx g0471(.A(n2276), .B(pi30), .O(n570));
  andx g0472(.A(pi27), .B(n192), .O(n571));
  andx g0473(.A(n1160), .B(n2342), .O(n572));
  andx g0474(.A(pi30), .B(pi31), .O(n573));
  andx g0475(.A(n2274), .B(n2383), .O(n574));
  andx g0476(.A(n2588), .B(n2342), .O(n575));
  andx g0477(.A(n261), .B(pi27), .O(n576));
  andx g0478(.A(n1161), .B(n2433), .O(n577));
  andx g0479(.A(n1162), .B(pi28), .O(n578));
  andx g0480(.A(n1159), .B(n2474), .O(n579));
  andx g0481(.A(n1163), .B(pi25), .O(n580));
  andx g0482(.A(n1166), .B(n1165), .O(n581));
  andx g0483(.A(n1168), .B(n1167), .O(n582));
  andx g0484(.A(n1170), .B(n1169), .O(n583));
  andx g0485(.A(n1172), .B(n1171), .O(n584));
  andx g0486(.A(n1164), .B(n2284), .O(n585));
  andx g0487(.A(n262), .B(pi26), .O(n586));
  andx g0488(.A(n1047), .B(pi27), .O(n587));
  andx g0489(.A(n171), .B(n2342), .O(n588));
  andx g0490(.A(n1029), .B(n2436), .O(n589));
  andx g0491(.A(n1173), .B(pi28), .O(n590));
  andx g0492(.A(n2307), .B(pi30), .O(n591));
  andx g0493(.A(n2289), .B(n2342), .O(n592));
  andx g0494(.A(n265), .B(pi27), .O(n593));
  andx g0495(.A(pi27), .B(n191), .O(n594));
  andx g0496(.A(n233), .B(n2343), .O(n595));
  andx g0497(.A(n1175), .B(n2434), .O(n596));
  andx g0498(.A(n264), .B(pi28), .O(n597));
  andx g0499(.A(n1174), .B(n2474), .O(n598));
  andx g0500(.A(n1176), .B(pi25), .O(n599));
  andx g0501(.A(n1179), .B(n1178), .O(n600));
  andx g0502(.A(n1181), .B(n1180), .O(n601));
  andx g0503(.A(n1183), .B(n1182), .O(n602));
  andx g0504(.A(n1177), .B(n2287), .O(n603));
  andx g0505(.A(n266), .B(pi26), .O(n604));
  andx g0506(.A(n2574), .B(pi25), .O(n605));
  andx g0507(.A(n2522), .B(n2474), .O(n606));
  andx g0508(.A(pi25), .B(n191), .O(n607));
  andx g0509(.A(n197), .B(n2475), .O(n608));
  andx g0510(.A(n1184), .B(n2343), .O(n609));
  andx g0511(.A(n1185), .B(pi27), .O(n610));
  andx g0512(.A(n2572), .B(pi25), .O(n611));
  andx g0513(.A(n177), .B(n2475), .O(n612));
  andx g0514(.A(n269), .B(n2343), .O(n613));
  andx g0515(.A(n1187), .B(pi27), .O(n614));
  andx g0516(.A(n1186), .B(n2440), .O(n615));
  andx g0517(.A(n1188), .B(pi28), .O(n616));
  andx g0518(.A(n1191), .B(n1190), .O(n617));
  andx g0519(.A(n1193), .B(n1192), .O(n618));
  andx g0520(.A(n1032), .B(n2434), .O(n619));
  andx g0521(.A(n268), .B(pi28), .O(n620));
  andx g0522(.A(n1189), .B(n2633), .O(n621));
  andx g0523(.A(n1194), .B(pi26), .O(n622));
  andx g0524(.A(n1112), .B(n2343), .O(n623));
  andx g0525(.A(pi27), .B(n2258), .O(n624));
  andx g0526(.A(n2403), .B(n2266), .O(n625));
  andx g0527(.A(pi30), .B(n2312), .O(n626));
  andx g0528(.A(n2280), .B(n2344), .O(n627));
  andx g0529(.A(n1196), .B(pi27), .O(n628));
  andx g0530(.A(n1195), .B(n2437), .O(n629));
  andx g0531(.A(n1197), .B(pi28), .O(n630));
  andx g0532(.A(n2581), .B(n2344), .O(n631));
  andx g0533(.A(n2586), .B(pi27), .O(n632));
  andx g0534(.A(n214), .B(n2348), .O(n633));
  andx g0535(.A(n1028), .B(pi27), .O(n634));
  andx g0536(.A(n1199), .B(n2434), .O(n635));
  andx g0537(.A(n1200), .B(pi28), .O(n636));
  andx g0538(.A(n1198), .B(n2475), .O(n637));
  andx g0539(.A(n1201), .B(pi25), .O(n638));
  andx g0540(.A(n1204), .B(n1203), .O(n639));
  andx g0541(.A(n1206), .B(n1205), .O(n640));
  andx g0542(.A(n1208), .B(n1207), .O(n641));
  andx g0543(.A(n1202), .B(n2259), .O(n642));
  andx g0544(.A(n271), .B(pi26), .O(n643));
  andx g0545(.A(n2317), .B(pi27), .O(n644));
  andx g0546(.A(n2587), .B(n2344), .O(n645));
  andx g0547(.A(pi31), .B(n2384), .O(n646));
  andx g0548(.A(pi30), .B(n2281), .O(n647));
  andx g0549(.A(n2314), .B(n2344), .O(n648));
  andx g0550(.A(n274), .B(pi27), .O(n649));
  andx g0551(.A(n1209), .B(n2437), .O(n650));
  andx g0552(.A(n1210), .B(pi28), .O(n651));
  andx g0553(.A(n2315), .B(n2383), .O(n652));
  andx g0554(.A(pi30), .B(n2275), .O(n653));
  andx g0555(.A(n1025), .B(n2673), .O(n654));
  andx g0556(.A(n1212), .B(pi27), .O(n655));
  andx g0557(.A(n2528), .B(pi27), .O(n656));
  andx g0558(.A(n1213), .B(n2434), .O(n657));
  andx g0559(.A(n1214), .B(pi28), .O(n658));
  andx g0560(.A(n1211), .B(n2475), .O(n659));
  andx g0561(.A(n1215), .B(pi25), .O(n660));
  andx g0562(.A(n1218), .B(n1217), .O(n661));
  andx g0563(.A(n1220), .B(n1219), .O(n662));
  andx g0564(.A(n1216), .B(n2295), .O(n663));
  andx g0565(.A(n275), .B(pi26), .O(n664));
  andx g0566(.A(n2584), .B(n2673), .O(n665));
  andx g0567(.A(n2522), .B(pi27), .O(n666));
  andx g0568(.A(n246), .B(pi27), .O(n667));
  andx g0569(.A(n1221), .B(n2448), .O(n668));
  andx g0570(.A(n1222), .B(pi28), .O(n669));
  andx g0571(.A(pi30), .B(n2321), .O(n670));
  andx g0572(.A(pi29), .B(n2386), .O(n671));
  andx g0573(.A(n2402), .B(n2320), .O(n672));
  andx g0574(.A(n2290), .B(pi30), .O(n673));
  andx g0575(.A(n277), .B(n2345), .O(n674));
  andx g0576(.A(n1224), .B(pi27), .O(n675));
  andx g0577(.A(n1225), .B(n2435), .O(n676));
  andx g0578(.A(n1033), .B(pi28), .O(n677));
  andx g0579(.A(n1223), .B(n2476), .O(n678));
  andx g0580(.A(n1226), .B(pi25), .O(n679));
  andx g0581(.A(n1229), .B(n1228), .O(n680));
  andx g0582(.A(n1231), .B(n1230), .O(n681));
  andx g0583(.A(n1233), .B(n1232), .O(n682));
  andx g0584(.A(n1227), .B(n2286), .O(n683));
  andx g0585(.A(n278), .B(pi26), .O(n684));
  andx g0586(.A(pi30), .B(n2279), .O(n685));
  andx g0587(.A(n2290), .B(n2385), .O(n686));
  andx g0588(.A(n280), .B(n2345), .O(n687));
  andx g0589(.A(n180), .B(pi27), .O(n688));
  andx g0590(.A(pi31), .B(n2384), .O(n689));
  andx g0591(.A(pi30), .B(n2302), .O(n690));
  andx g0592(.A(n251), .B(pi27), .O(n691));
  andx g0593(.A(n1235), .B(n2345), .O(n692));
  andx g0594(.A(n1234), .B(n2438), .O(n693));
  andx g0595(.A(n1236), .B(pi28), .O(n694));
  andx g0596(.A(n2530), .B(n2345), .O(n695));
  andx g0597(.A(n2538), .B(pi27), .O(n696));
  orx  g0598(.A(n2282), .B(n2405), .O(n697));
  andx g0599(.A(n2559), .B(pi27), .O(n698));
  andx g0600(.A(n211), .B(n2346), .O(n699));
  andx g0601(.A(n1238), .B(n2441), .O(n700));
  andx g0602(.A(n1239), .B(pi28), .O(n701));
  andx g0603(.A(n1237), .B(n2476), .O(n702));
  andx g0604(.A(n1240), .B(pi25), .O(n703));
  andx g0605(.A(n1243), .B(n1242), .O(n704));
  andx g0606(.A(n1245), .B(n1244), .O(n705));
  andx g0607(.A(n1247), .B(n1246), .O(n706));
  andx g0608(.A(n1241), .B(n2259), .O(n707));
  andx g0609(.A(n281), .B(pi26), .O(n708));
  andx g0610(.A(n2303), .B(n2476), .O(n709));
  andx g0611(.A(pi25), .B(n198), .O(n710));
  andx g0612(.A(pi30), .B(n2320), .O(n711));
  andx g0613(.A(n2312), .B(n2384), .O(n712));
  andx g0614(.A(n227), .B(pi25), .O(n713));
  andx g0615(.A(n284), .B(n2476), .O(n714));
  andx g0616(.A(n1248), .B(n2346), .O(n715));
  andx g0617(.A(n1249), .B(pi27), .O(n716));
  andx g0618(.A(n211), .B(pi25), .O(n717));
  andx g0619(.A(n194), .B(n2477), .O(n718));
  andx g0620(.A(n2584), .B(pi27), .O(n719));
  andx g0621(.A(n1251), .B(n2346), .O(n720));
  andx g0622(.A(n1250), .B(n2438), .O(n721));
  andx g0623(.A(n1252), .B(pi28), .O(n722));
  andx g0624(.A(pi30), .B(n2293), .O(n723));
  andx g0625(.A(n2313), .B(n2385), .O(n724));
  andx g0626(.A(n1255), .B(n1254), .O(n725));
  andx g0627(.A(n1257), .B(n1256), .O(n726));
  andx g0628(.A(n1253), .B(n2262), .O(n727));
  andx g0629(.A(n285), .B(pi26), .O(n728));
  andx g0630(.A(n2613), .B(n2346), .O(n729));
  andx g0631(.A(pi27), .B(n2531), .O(n730));
  andx g0632(.A(n1258), .B(n2443), .O(n731));
  andx g0633(.A(n290), .B(pi28), .O(n732));
  orx  g0634(.A(n2546), .B(n2357), .O(n733));
  andx g0635(.A(n1261), .B(n1260), .O(n734));
  andx g0636(.A(n2277), .B(pi30), .O(n735));
  andx g0637(.A(n2313), .B(n2385), .O(n736));
  andx g0638(.A(n1263), .B(n1262), .O(n737));
  andx g0639(.A(n1259), .B(n2477), .O(n738));
  andx g0640(.A(n291), .B(pi25), .O(n739));
  andx g0641(.A(n2281), .B(n2385), .O(n740));
  andx g0642(.A(n1266), .B(n1265), .O(n741));
  andx g0643(.A(n1268), .B(n1267), .O(n742));
  andx g0644(.A(n1270), .B(n1269), .O(n743));
  andx g0645(.A(n1264), .B(n2259), .O(n744));
  andx g0646(.A(n292), .B(pi26), .O(n745));
  andx g0647(.A(pi30), .B(pi31), .O(n746));
  andx g0648(.A(n2302), .B(n2387), .O(n747));
  andx g0649(.A(n1072), .B(pi25), .O(n748));
  andx g0650(.A(n1271), .B(n2477), .O(n749));
  andx g0651(.A(n2525), .B(n2477), .O(n750));
  andx g0652(.A(n2540), .B(pi25), .O(n751));
  andx g0653(.A(n1272), .B(n2349), .O(n752));
  andx g0654(.A(n1273), .B(pi27), .O(n753));
  andx g0655(.A(n242), .B(pi25), .O(n754));
  andx g0656(.A(n2567), .B(n2478), .O(n755));
  andx g0657(.A(pi25), .B(n196), .O(n756));
  andx g0658(.A(n1165), .B(n2478), .O(n757));
  andx g0659(.A(n1275), .B(n2347), .O(n758));
  andx g0660(.A(n1276), .B(pi27), .O(n759));
  andx g0661(.A(n1274), .B(n2435), .O(n760));
  andx g0662(.A(n1277), .B(pi28), .O(n761));
  andx g0663(.A(n1280), .B(n1279), .O(n762));
  andx g0664(.A(n1282), .B(n1281), .O(n763));
  andx g0665(.A(n1278), .B(n2285), .O(n764));
  andx g0666(.A(n294), .B(pi26), .O(n765));
  andx g0667(.A(n265), .B(pi25), .O(n766));
  andx g0668(.A(n1037), .B(n2478), .O(n767));
  andx g0669(.A(pi30), .B(pi31), .O(n768));
  andx g0670(.A(n2312), .B(n2386), .O(n769));
  andx g0671(.A(n2577), .B(n2478), .O(n770));
  andx g0672(.A(n297), .B(pi25), .O(n771));
  andx g0673(.A(n1283), .B(n2355), .O(n772));
  andx g0674(.A(n1284), .B(pi27), .O(n773));
  andx g0675(.A(n2280), .B(n2386), .O(n774));
  andx g0676(.A(pi30), .B(n2274), .O(n775));
  andx g0677(.A(n251), .B(pi25), .O(n776));
  andx g0678(.A(n296), .B(n2479), .O(n777));
  andx g0679(.A(pi31), .B(n2387), .O(n778));
  andx g0680(.A(n2289), .B(pi30), .O(n779));
  andx g0681(.A(n288), .B(pi25), .O(n780));
  andx g0682(.A(n1287), .B(n2479), .O(n781));
  andx g0683(.A(n1286), .B(n2340), .O(n782));
  andx g0684(.A(n1288), .B(pi27), .O(n783));
  andx g0685(.A(n1285), .B(n2668), .O(n784));
  andx g0686(.A(n1289), .B(pi28), .O(n785));
  andx g0687(.A(n1292), .B(n1291), .O(n786));
  andx g0688(.A(n1294), .B(n1293), .O(n787));
  andx g0689(.A(n1296), .B(n1295), .O(n788));
  andx g0690(.A(n1290), .B(n2259), .O(n789));
  andx g0691(.A(n298), .B(pi26), .O(n790));
  andx g0692(.A(n2555), .B(n2479), .O(n791));
  andx g0693(.A(n2554), .B(pi25), .O(n792));
  andx g0694(.A(n1299), .B(n1298), .O(n793));
  andx g0695(.A(n2544), .B(n2479), .O(n794));
  andx g0696(.A(n793), .B(pi25), .O(n795));
  andx g0697(.A(n1297), .B(n2347), .O(n796));
  andx g0698(.A(n1300), .B(pi27), .O(n797));
  andx g0699(.A(pi30), .B(n2292), .O(n798));
  andx g0700(.A(n2317), .B(n2386), .O(n799));
  andx g0701(.A(n1031), .B(n2480), .O(n800));
  andx g0702(.A(n301), .B(pi25), .O(n801));
  andx g0703(.A(pi30), .B(n2315), .O(n802));
  andx g0704(.A(n2303), .B(n2387), .O(n803));
  andx g0705(.A(n202), .B(n2480), .O(n804));
  andx g0706(.A(n2551), .B(pi25), .O(n805));
  andx g0707(.A(n1302), .B(n2347), .O(n806));
  andx g0708(.A(n1303), .B(pi27), .O(n807));
  andx g0709(.A(n1301), .B(n2439), .O(n808));
  andx g0710(.A(n1304), .B(pi28), .O(n809));
  andx g0711(.A(n1307), .B(n1306), .O(n810));
  andx g0712(.A(n1309), .B(n1308), .O(n811));
  andx g0713(.A(n1311), .B(n1310), .O(n812));
  andx g0714(.A(n1305), .B(n2633), .O(n813));
  andx g0715(.A(n302), .B(pi26), .O(n814));
  andx g0716(.A(n2575), .B(pi27), .O(n815));
  andx g0717(.A(n200), .B(n2347), .O(n816));
  andx g0718(.A(pi27), .B(pi31), .O(n817));
  andx g0719(.A(n2576), .B(n2347), .O(n818));
  andx g0720(.A(n1312), .B(n2436), .O(n819));
  andx g0721(.A(n1313), .B(pi28), .O(n820));
  andx g0722(.A(pi31), .B(n2387), .O(n821));
  andx g0723(.A(n166), .B(pi30), .O(n822));
  andx g0724(.A(pi27), .B(n2318), .O(n823));
  andx g0725(.A(n1315), .B(n2348), .O(n824));
  andx g0726(.A(n261), .B(n2348), .O(n825));
  andx g0727(.A(n1212), .B(pi27), .O(n826));
  andx g0728(.A(n1316), .B(n2436), .O(n827));
  andx g0729(.A(n1317), .B(pi28), .O(n828));
  andx g0730(.A(n1314), .B(n2480), .O(n829));
  andx g0731(.A(n1318), .B(pi25), .O(n830));
  andx g0732(.A(n1321), .B(n1320), .O(n831));
  andx g0733(.A(n1323), .B(n1322), .O(n832));
  andx g0734(.A(n1325), .B(n1324), .O(n833));
  andx g0735(.A(n1327), .B(n1326), .O(n834));
  andx g0736(.A(n1319), .B(n2286), .O(n835));
  andx g0737(.A(n304), .B(pi26), .O(n836));
  andx g0738(.A(n2568), .B(pi28), .O(n837));
  andx g0739(.A(n2556), .B(n2451), .O(n838));
  andx g0740(.A(n1329), .B(n1328), .O(n839));
  andx g0741(.A(n173), .B(n2348), .O(n840));
  andx g0742(.A(pi27), .B(n203), .O(n841));
  andx g0743(.A(n213), .B(n2349), .O(n842));
  andx g0744(.A(n2558), .B(pi27), .O(n843));
  andx g0745(.A(n1330), .B(n2437), .O(n844));
  andx g0746(.A(n1331), .B(pi28), .O(n845));
  andx g0747(.A(n307), .B(n2480), .O(n846));
  andx g0748(.A(n1332), .B(pi25), .O(n847));
  andx g0749(.A(n1335), .B(n1334), .O(n848));
  andx g0750(.A(n1337), .B(n2258), .O(n849));
  andx g0751(.A(n1339), .B(n1338), .O(n850));
  andx g0752(.A(n1341), .B(n1340), .O(n851));
  andx g0753(.A(n1333), .B(n2287), .O(n852));
  andx g0754(.A(n308), .B(pi26), .O(n853));
  andx g0755(.A(n2577), .B(pi25), .O(n854));
  andx g0756(.A(n2624), .B(n2481), .O(n855));
  andx g0757(.A(n1039), .B(n2349), .O(n856));
  andx g0758(.A(n1342), .B(pi27), .O(n857));
  andx g0759(.A(n236), .B(pi25), .O(n858));
  andx g0760(.A(n204), .B(n2481), .O(n859));
  andx g0761(.A(n2522), .B(n2481), .O(n860));
  andx g0762(.A(n2585), .B(pi25), .O(n861));
  andx g0763(.A(n1344), .B(n2349), .O(n862));
  andx g0764(.A(n1345), .B(pi27), .O(n863));
  andx g0765(.A(n1343), .B(n2440), .O(n864));
  andx g0766(.A(n1346), .B(pi28), .O(n865));
  andx g0767(.A(n1349), .B(n1348), .O(n866));
  andx g0768(.A(n1351), .B(n1350), .O(n867));
  andx g0769(.A(n1353), .B(n1352), .O(n868));
  andx g0770(.A(n1347), .B(n2294), .O(n869));
  andx g0771(.A(n310), .B(pi26), .O(n870));
  andx g0772(.A(n207), .B(n2349), .O(n871));
  andx g0773(.A(n1315), .B(pi27), .O(n872));
  andx g0774(.A(n257), .B(pi27), .O(n873));
  andx g0775(.A(n2552), .B(n2350), .O(n874));
  andx g0776(.A(n1354), .B(n2437), .O(n875));
  andx g0777(.A(n1355), .B(pi28), .O(n876));
  andx g0778(.A(pi30), .B(pi31), .O(n877));
  andx g0779(.A(n205), .B(n2388), .O(n878));
  orx  g0780(.A(n2376), .B(n2274), .O(n879));
  andx g0781(.A(n2549), .B(pi27), .O(n880));
  andx g0782(.A(n313), .B(n2350), .O(n881));
  andx g0783(.A(n1040), .B(n2440), .O(n882));
  andx g0784(.A(n1357), .B(pi28), .O(n883));
  andx g0785(.A(n1356), .B(n2481), .O(n884));
  andx g0786(.A(n1358), .B(pi25), .O(n885));
  andx g0787(.A(n1361), .B(n1360), .O(n886));
  andx g0788(.A(n1359), .B(n2633), .O(n887));
  andx g0789(.A(n314), .B(pi26), .O(n888));
  andx g0790(.A(pi30), .B(n2282), .O(n889));
  andx g0791(.A(n2302), .B(n2388), .O(n890));
  andx g0792(.A(pi27), .B(n2516), .O(n891));
  andx g0793(.A(n318), .B(n2350), .O(n892));
  andx g0794(.A(n1362), .B(n2438), .O(n893));
  andx g0795(.A(n319), .B(pi28), .O(n894));
  orx  g0796(.A(pi30), .B(n2281), .O(n895));
  andx g0797(.A(n164), .B(n2350), .O(n896));
  andx g0798(.A(n2521), .B(pi27), .O(n897));
  andx g0799(.A(pi30), .B(n2303), .O(n898));
  andx g0800(.A(n2316), .B(n2388), .O(n899));
  andx g0801(.A(n173), .B(pi27), .O(n900));
  andx g0802(.A(n317), .B(n2351), .O(n901));
  andx g0803(.A(n1364), .B(n2440), .O(n902));
  andx g0804(.A(n1365), .B(pi28), .O(n903));
  andx g0805(.A(n1363), .B(n2482), .O(n904));
  andx g0806(.A(n1366), .B(pi25), .O(n905));
  orx  g0807(.A(n2528), .B(n2357), .O(n906));
  andx g0808(.A(n1369), .B(n1368), .O(n907));
  andx g0809(.A(n1367), .B(n2261), .O(n908));
  andx g0810(.A(n320), .B(pi26), .O(n909));
  andx g0811(.A(n1235), .B(n2351), .O(n910));
  andx g0812(.A(n2547), .B(pi27), .O(n911));
  andx g0813(.A(n2603), .B(pi27), .O(n912));
  andx g0814(.A(n235), .B(n2351), .O(n913));
  andx g0815(.A(n1370), .B(n2439), .O(n914));
  andx g0816(.A(n1371), .B(pi28), .O(n915));
  andx g0817(.A(n2524), .B(pi27), .O(n916));
  andx g0818(.A(n1037), .B(n2352), .O(n917));
  andx g0819(.A(n2582), .B(pi27), .O(n918));
  andx g0820(.A(n1042), .B(n2351), .O(n919));
  andx g0821(.A(n1373), .B(n2439), .O(n920));
  andx g0822(.A(n1374), .B(pi28), .O(n921));
  andx g0823(.A(n1372), .B(n2482), .O(n922));
  andx g0824(.A(n1375), .B(pi25), .O(n923));
  andx g0825(.A(n1378), .B(n1377), .O(n924));
  andx g0826(.A(n1380), .B(n1379), .O(n925));
  andx g0827(.A(n1382), .B(n1381), .O(n926));
  andx g0828(.A(n1376), .B(n2286), .O(n927));
  andx g0829(.A(n322), .B(pi26), .O(n928));
  andx g0830(.A(n206), .B(n2352), .O(n929));
  andx g0831(.A(pi27), .B(n199), .O(n930));
  andx g0832(.A(n1043), .B(n2442), .O(n931));
  andx g0833(.A(n1383), .B(pi28), .O(n932));
  andx g0834(.A(n2532), .B(n2352), .O(n933));
  andx g0835(.A(n265), .B(pi27), .O(n934));
  andx g0836(.A(n1385), .B(n2434), .O(n935));
  andx g0837(.A(n1044), .B(pi28), .O(n936));
  andx g0838(.A(n1384), .B(n2482), .O(n937));
  andx g0839(.A(n1386), .B(pi25), .O(n938));
  andx g0840(.A(n1389), .B(n1388), .O(n939));
  andx g0841(.A(n1391), .B(n1390), .O(n940));
  andx g0842(.A(n1393), .B(n1392), .O(n941));
  andx g0843(.A(n1387), .B(n2284), .O(n942));
  andx g0844(.A(n324), .B(pi26), .O(n943));
  andx g0845(.A(n2545), .B(n2353), .O(n944));
  andx g0846(.A(n2565), .B(pi27), .O(n945));
  andx g0847(.A(n2603), .B(n2353), .O(n946));
  andx g0848(.A(n2548), .B(pi27), .O(n947));
  andx g0849(.A(n1394), .B(n2441), .O(n948));
  andx g0850(.A(n1395), .B(pi28), .O(n949));
  andx g0851(.A(n2584), .B(n2352), .O(n950));
  andx g0852(.A(n2557), .B(pi27), .O(n951));
  andx g0853(.A(n2551), .B(n2353), .O(n952));
  andx g0854(.A(n2550), .B(pi27), .O(n953));
  andx g0855(.A(n1397), .B(n2441), .O(n954));
  andx g0856(.A(n1398), .B(pi28), .O(n955));
  andx g0857(.A(n1396), .B(n2483), .O(n956));
  andx g0858(.A(n1399), .B(pi25), .O(n957));
  andx g0859(.A(n1402), .B(n1401), .O(n958));
  andx g0860(.A(n1404), .B(n1403), .O(n959));
  andx g0861(.A(n1400), .B(n2260), .O(n960));
  andx g0862(.A(n327), .B(pi26), .O(n961));
  andx g0863(.A(pi29), .B(n2388), .O(n962));
  andx g0864(.A(pi30), .B(n1972), .O(n963));
  andx g0865(.A(n2569), .B(pi28), .O(n964));
  andx g0866(.A(n1405), .B(n2441), .O(n965));
  andx g0867(.A(n2582), .B(pi28), .O(n966));
  andx g0868(.A(n2588), .B(n2442), .O(n967));
  andx g0869(.A(n1406), .B(n2354), .O(n968));
  andx g0870(.A(n1407), .B(pi27), .O(n969));
  andx g0871(.A(n195), .B(n2442), .O(n970));
  andx g0872(.A(n2554), .B(pi28), .O(n971));
  andx g0873(.A(pi27), .B(n2258), .O(n972));
  andx g0874(.A(n1409), .B(n2354), .O(n973));
  andx g0875(.A(n1408), .B(n2483), .O(n974));
  andx g0876(.A(n1410), .B(pi25), .O(n975));
  andx g0877(.A(n1413), .B(n1412), .O(n976));
  andx g0878(.A(n1415), .B(n1414), .O(n977));
  andx g0879(.A(n1411), .B(n2261), .O(n978));
  andx g0880(.A(n330), .B(pi26), .O(n979));
  andx g0881(.A(n2581), .B(pi26), .O(n980));
  andx g0882(.A(n2563), .B(n2285), .O(n981));
  andx g0883(.A(n1046), .B(n2354), .O(n982));
  andx g0884(.A(n1416), .B(pi27), .O(n983));
  andx g0885(.A(n2583), .B(n2261), .O(n984));
  andx g0886(.A(n1196), .B(pi26), .O(n985));
  andx g0887(.A(n2283), .B(n2262), .O(n986));
  andx g0888(.A(pi26), .B(n2532), .O(n987));
  andx g0889(.A(n1418), .B(n2355), .O(n988));
  andx g0890(.A(n1419), .B(pi27), .O(n989));
  andx g0891(.A(n1417), .B(n2442), .O(n990));
  andx g0892(.A(n1420), .B(pi28), .O(n991));
  andx g0893(.A(n1423), .B(n1422), .O(n992));
  andx g0894(.A(n1425), .B(n1424), .O(n993));
  andx g0895(.A(n1427), .B(n1426), .O(n994));
  andx g0896(.A(n1421), .B(n2483), .O(n995));
  andx g0897(.A(n332), .B(pi25), .O(n996));
  andx g0898(.A(n233), .B(n2284), .O(n997));
  andx g0899(.A(n1224), .B(pi26), .O(n998));
  andx g0900(.A(n2582), .B(n2287), .O(n999));
  andx g0901(.A(pi26), .B(n2258), .O(n1000));
  andx g0902(.A(n1428), .B(n2355), .O(n1001));
  andx g0903(.A(n1429), .B(pi27), .O(n1002));
  andx g0904(.A(n2313), .B(n2294), .O(n1003));
  andx g0905(.A(n1112), .B(pi26), .O(n1004));
  andx g0906(.A(n2525), .B(pi26), .O(n1005));
  andx g0907(.A(n2566), .B(n2261), .O(n1006));
  andx g0908(.A(n1431), .B(n2355), .O(n1007));
  andx g0909(.A(n1432), .B(pi27), .O(n1008));
  andx g0910(.A(n1430), .B(n2443), .O(n1009));
  andx g0911(.A(n1433), .B(pi28), .O(n1010));
  andx g0912(.A(n1436), .B(n1435), .O(n1011));
  andx g0913(.A(n1438), .B(n1437), .O(n1012));
  andx g0914(.A(n1434), .B(n2483), .O(n1013));
  andx g0915(.A(n334), .B(pi25), .O(n1014));
  orx  g0916(.A(pi29), .B(pi30), .O(n1015));
  orx  g0917(.A(pi27), .B(n2283), .O(n1016));
  orx  g0918(.A(n2523), .B(n2357), .O(n1017));
  orx  g0919(.A(n2525), .B(n2359), .O(n1018));
  orx  g0920(.A(n2317), .B(n2404), .O(n1019));
  orx  g0921(.A(n343), .B(n189), .O(n1020));
  orx  g0922(.A(n2549), .B(n165), .O(n1021));
  orx  g0923(.A(n2593), .B(n168), .O(n1022));
  orx  g0924(.A(n2521), .B(n2287), .O(n1023));
  orx  g0925(.A(n2289), .B(n2404), .O(n1024));
  orx  g0926(.A(n2276), .B(n2405), .O(n1025));
  orx  g0927(.A(n172), .B(n2573), .O(n1026));
  orx  g0928(.A(n2521), .B(n2358), .O(n1027));
  orx  g0929(.A(n2275), .B(pi30), .O(n1028));
  orx  g0930(.A(n175), .B(n2572), .O(n1029));
  orx  g0931(.A(n176), .B(n2497), .O(n1030));
  orx  g0932(.A(n2307), .B(n2404), .O(n1031));
  orx  g0933(.A(n179), .B(n178), .O(n1032));
  orx  g0934(.A(n2526), .B(n209), .O(n1033));
  orx  g0935(.A(n182), .B(n181), .O(n1034));
  orx  g0936(.A(n207), .B(n2357), .O(n1035));
  orx  g0937(.A(n183), .B(n181), .O(n1036));
  orx  g0938(.A(n2613), .B(n2276), .O(n1037));
  orx  g0939(.A(n2334), .B(n306), .O(n1038));
  orx  g0940(.A(n184), .B(n2528), .O(n1039));
  orx  g0941(.A(n185), .B(n2521), .O(n1040));
  orx  g0942(.A(n265), .B(n2358), .O(n1041));
  orx  g0943(.A(n2559), .B(n2308), .O(n1042));
  orx  g0944(.A(n186), .B(n2546), .O(n1043));
  orx  g0945(.A(n187), .B(n2549), .O(n1044));
  orx  g0946(.A(n2521), .B(n2454), .O(n1045));
  orx  g0947(.A(n188), .B(n2521), .O(n1046));
  orx  g0948(.A(n350), .B(n351), .O(n1047));
  orx  g0949(.A(n352), .B(n353), .O(n1048));
  orx  g0950(.A(n354), .B(n355), .O(n1049));
  orx  g0951(.A(n356), .B(n357), .O(n1050));
  orx  g0952(.A(n360), .B(n361), .O(n1051));
  orx  g0953(.A(n362), .B(n363), .O(n1052));
  orx  g0954(.A(n364), .B(n365), .O(n1053));
  orx  g0955(.A(pi27), .B(n212), .O(n1054));
  orx  g0956(.A(n2330), .B(n211), .O(n1055));
  orx  g0957(.A(pi28), .B(n369), .O(n1056));
  orx  g0958(.A(n2418), .B(n210), .O(n1057));
  orx  g0959(.A(n379), .B(n380), .O(n1058));
  orx  g0960(.A(n381), .B(n382), .O(n1059));
  orx  g0961(.A(n383), .B(n384), .O(n1060));
  orx  g0962(.A(n385), .B(n386), .O(n1061));
  orx  g0963(.A(n387), .B(n388), .O(n1062));
  orx  g0964(.A(n389), .B(n390), .O(n1063));
  orx  g0965(.A(pi27), .B(n219), .O(n1064));
  orx  g0966(.A(n2334), .B(n218), .O(n1065));
  orx  g0967(.A(pi27), .B(n209), .O(n1066));
  orx  g0968(.A(n2530), .B(n2357), .O(n1067));
  orx  g0969(.A(pi28), .B(n395), .O(n1068));
  orx  g0970(.A(n2418), .B(n396), .O(n1069));
  orx  g0971(.A(pi31), .B(n2404), .O(n1070));
  orx  g0972(.A(pi30), .B(n2283), .O(n1071));
  orx  g0973(.A(n401), .B(n402), .O(n1072));
  orx  g0974(.A(n404), .B(n403), .O(n1073));
  orx  g0975(.A(n405), .B(n406), .O(n1074));
  orx  g0976(.A(n407), .B(n408), .O(n1075));
  orx  g0977(.A(n410), .B(n409), .O(n1076));
  orx  g0978(.A(n411), .B(n412), .O(n1077));
  orx  g0979(.A(n413), .B(n414), .O(n1078));
  orx  g0980(.A(pi31), .B(n2405), .O(n1079));
  orx  g0981(.A(pi30), .B(n2280), .O(n1080));
  orx  g0982(.A(pi27), .B(n415), .O(n1081));
  orx  g0983(.A(n2520), .B(n2356), .O(n1082));
  orx  g0984(.A(pi31), .B(pi27), .O(n1083));
  orx  g0985(.A(n2589), .B(n2358), .O(n1084));
  orx  g0986(.A(pi28), .B(n416), .O(n1085));
  orx  g0987(.A(n2418), .B(n417), .O(n1086));
  orx  g0988(.A(n421), .B(n422), .O(n1087));
  orx  g0989(.A(n423), .B(n424), .O(n1088));
  orx  g0990(.A(n427), .B(n428), .O(n1089));
  orx  g0991(.A(n431), .B(n432), .O(n1090));
  orx  g0992(.A(n433), .B(n434), .O(n1091));
  orx  g0993(.A(n435), .B(n436), .O(n1092));
  orx  g0994(.A(pi27), .B(n228), .O(n1093));
  orx  g0995(.A(n2334), .B(n227), .O(n1094));
  orx  g0996(.A(pi27), .B(n2530), .O(n1095));
  orx  g0997(.A(n2525), .B(n2359), .O(n1096));
  orx  g0998(.A(pi28), .B(n441), .O(n1097));
  orx  g0999(.A(n2419), .B(n442), .O(n1098));
  orx  g1000(.A(n449), .B(n450), .O(n1099));
  orx  g1001(.A(n453), .B(n454), .O(n1100));
  orx  g1002(.A(n455), .B(n456), .O(n1101));
  orx  g1003(.A(n459), .B(n460), .O(n1102));
  orx  g1004(.A(n461), .B(n462), .O(n1103));
  orx  g1005(.A(n463), .B(n464), .O(n1104));
  orx  g1006(.A(n465), .B(n466), .O(n1105));
  orx  g1007(.A(pi27), .B(n235), .O(n1106));
  orx  g1008(.A(n2333), .B(n234), .O(n1107));
  orx  g1009(.A(n2520), .B(n2358), .O(n1108));
  orx  g1010(.A(pi27), .B(n233), .O(n1109));
  orx  g1011(.A(pi28), .B(n471), .O(n1110));
  orx  g1012(.A(n2419), .B(n474), .O(n1111));
  orx  g1013(.A(n478), .B(n479), .O(n1112));
  orx  g1014(.A(n482), .B(n483), .O(n1113));
  orx  g1015(.A(n486), .B(n487), .O(n1114));
  orx  g1016(.A(n488), .B(n489), .O(n1115));
  orx  g1017(.A(n490), .B(n491), .O(n1116));
  orx  g1018(.A(n494), .B(n495), .O(n1117));
  orx  g1019(.A(n496), .B(n497), .O(n1118));
  orx  g1020(.A(n498), .B(n499), .O(n1119));
  orx  g1021(.A(pi27), .B(n2276), .O(n1120));
  orx  g1022(.A(n2333), .B(n2582), .O(n1121));
  orx  g1023(.A(n2419), .B(n210), .O(n1122));
  orx  g1024(.A(pi28), .B(n500), .O(n1123));
  orx  g1025(.A(n504), .B(n505), .O(n1124));
  orx  g1026(.A(n506), .B(n507), .O(n1125));
  orx  g1027(.A(n625), .B(n508), .O(n1126));
  orx  g1028(.A(n511), .B(n512), .O(n1127));
  orx  g1029(.A(n513), .B(n514), .O(n1128));
  orx  g1030(.A(n515), .B(n516), .O(n1129));
  orx  g1031(.A(pi28), .B(n2569), .O(n1130));
  orx  g1032(.A(n2522), .B(n2455), .O(n1131));
  orx  g1033(.A(n2528), .B(n2452), .O(n1132));
  orx  g1034(.A(pi28), .B(n246), .O(n1133));
  orx  g1035(.A(pi27), .B(n517), .O(n1134));
  orx  g1036(.A(n2333), .B(n520), .O(n1135));
  orx  g1037(.A(n526), .B(n527), .O(n1136));
  orx  g1038(.A(n528), .B(n529), .O(n1137));
  orx  g1039(.A(n530), .B(n531), .O(n1138));
  orx  g1040(.A(n534), .B(n535), .O(n1139));
  orx  g1041(.A(n536), .B(n537), .O(n1140));
  orx  g1042(.A(n538), .B(n539), .O(n1141));
  orx  g1043(.A(pi28), .B(n542), .O(n1142));
  orx  g1044(.A(n2419), .B(n250), .O(n1143));
  orx  g1045(.A(n547), .B(n548), .O(n1144));
  orx  g1046(.A(n549), .B(n550), .O(n1145));
  orx  g1047(.A(pi30), .B(n2266), .O(n1146));
  orx  g1048(.A(pi29), .B(n2404), .O(n1147));
  orx  g1049(.A(n552), .B(n553), .O(n1148));
  orx  g1050(.A(n555), .B(n556), .O(n1149));
  orx  g1051(.A(n557), .B(n558), .O(n1150));
  orx  g1052(.A(n559), .B(n560), .O(n1151));
  orx  g1053(.A(n2333), .B(n2532), .O(n1152));
  orx  g1054(.A(pi27), .B(n2567), .O(n1153));
  orx  g1055(.A(pi28), .B(n561), .O(n1154));
  orx  g1056(.A(n2420), .B(n256), .O(n1155));
  orx  g1057(.A(n565), .B(n535), .O(n1156));
  orx  g1058(.A(n2326), .B(n242), .O(n1157));
  orx  g1059(.A(pi27), .B(n2570), .O(n1158));
  orx  g1060(.A(n567), .B(n568), .O(n1159));
  orx  g1061(.A(n569), .B(n570), .O(n1160));
  orx  g1062(.A(n571), .B(n572), .O(n1161));
  orx  g1063(.A(n575), .B(n576), .O(n1162));
  orx  g1064(.A(n577), .B(n578), .O(n1163));
  orx  g1065(.A(n579), .B(n580), .O(n1164));
  orx  g1066(.A(n2279), .B(n2403), .O(n1165));
  orx  g1067(.A(pi30), .B(n2275), .O(n1166));
  orx  g1068(.A(pi27), .B(n242), .O(n1167));
  orx  g1069(.A(n2332), .B(n581), .O(n1168));
  orx  g1070(.A(n2520), .B(n2345), .O(n1169));
  orx  g1071(.A(pi27), .B(n2257), .O(n1170));
  orx  g1072(.A(pi28), .B(n582), .O(n1171));
  orx  g1073(.A(n2420), .B(n583), .O(n1172));
  orx  g1074(.A(n587), .B(n588), .O(n1173));
  orx  g1075(.A(n589), .B(n590), .O(n1174));
  orx  g1076(.A(n592), .B(n593), .O(n1175));
  orx  g1077(.A(n596), .B(n597), .O(n1176));
  orx  g1078(.A(n598), .B(n599), .O(n1177));
  orx  g1079(.A(pi27), .B(n2579), .O(n1178));
  orx  g1080(.A(n2332), .B(n233), .O(n1179));
  orx  g1081(.A(n2525), .B(n2360), .O(n1180));
  orx  g1082(.A(pi27), .B(n239), .O(n1181));
  orx  g1083(.A(pi28), .B(n600), .O(n1182));
  orx  g1084(.A(n2420), .B(n601), .O(n1183));
  orx  g1085(.A(n605), .B(n606), .O(n1184));
  orx  g1086(.A(n607), .B(n608), .O(n1185));
  orx  g1087(.A(n609), .B(n610), .O(n1186));
  orx  g1088(.A(n611), .B(n612), .O(n1187));
  orx  g1089(.A(n613), .B(n614), .O(n1188));
  orx  g1090(.A(n615), .B(n616), .O(n1189));
  orx  g1091(.A(n2320), .B(n2405), .O(n1190));
  orx  g1092(.A(pi30), .B(n2302), .O(n1191));
  orx  g1093(.A(pi27), .B(n2585), .O(n1192));
  orx  g1094(.A(n2524), .B(n2359), .O(n1193));
  orx  g1095(.A(n619), .B(n620), .O(n1194));
  orx  g1096(.A(n623), .B(n624), .O(n1195));
  orx  g1097(.A(n625), .B(n626), .O(n1196));
  orx  g1098(.A(n627), .B(n628), .O(n1197));
  orx  g1099(.A(n629), .B(n630), .O(n1198));
  orx  g1100(.A(n631), .B(n632), .O(n1199));
  orx  g1101(.A(n633), .B(n634), .O(n1200));
  orx  g1102(.A(n635), .B(n636), .O(n1201));
  orx  g1103(.A(n637), .B(n638), .O(n1202));
  orx  g1104(.A(n2332), .B(n212), .O(n1203));
  orx  g1105(.A(pi27), .B(n2545), .O(n1204));
  orx  g1106(.A(n2530), .B(n2359), .O(n1205));
  orx  g1107(.A(pi27), .B(n257), .O(n1206));
  orx  g1108(.A(pi28), .B(n639), .O(n1207));
  orx  g1109(.A(n2420), .B(n640), .O(n1208));
  orx  g1110(.A(n644), .B(n645), .O(n1209));
  orx  g1111(.A(n648), .B(n649), .O(n1210));
  orx  g1112(.A(n650), .B(n651), .O(n1211));
  orx  g1113(.A(n652), .B(n653), .O(n1212));
  orx  g1114(.A(n654), .B(n655), .O(n1213));
  orx  g1115(.A(n386), .B(n656), .O(n1214));
  orx  g1116(.A(n657), .B(n658), .O(n1215));
  orx  g1117(.A(n659), .B(n660), .O(n1216));
  orx  g1118(.A(n2329), .B(n2564), .O(n1217));
  orx  g1119(.A(pi27), .B(n273), .O(n1218));
  orx  g1120(.A(n2421), .B(n250), .O(n1219));
  orx  g1121(.A(pi28), .B(n661), .O(n1220));
  orx  g1122(.A(n665), .B(n666), .O(n1221));
  orx  g1123(.A(n1612), .B(n667), .O(n1222));
  orx  g1124(.A(n668), .B(n669), .O(n1223));
  orx  g1125(.A(n672), .B(n673), .O(n1224));
  orx  g1126(.A(n674), .B(n675), .O(n1225));
  orx  g1127(.A(n676), .B(n677), .O(n1226));
  orx  g1128(.A(n678), .B(n679), .O(n1227));
  orx  g1129(.A(pi27), .B(n169), .O(n1228));
  orx  g1130(.A(n2332), .B(n219), .O(n1229));
  orx  g1131(.A(n2330), .B(n2532), .O(n1230));
  orx  g1132(.A(pi27), .B(n257), .O(n1231));
  orx  g1133(.A(pi28), .B(n680), .O(n1232));
  orx  g1134(.A(n2421), .B(n681), .O(n1233));
  orx  g1135(.A(n687), .B(n688), .O(n1234));
  orx  g1136(.A(n689), .B(n690), .O(n1235));
  orx  g1137(.A(n691), .B(n692), .O(n1236));
  orx  g1138(.A(n693), .B(n694), .O(n1237));
  orx  g1139(.A(n695), .B(n696), .O(n1238));
  orx  g1140(.A(n698), .B(n699), .O(n1239));
  orx  g1141(.A(n700), .B(n701), .O(n1240));
  orx  g1142(.A(n702), .B(n703), .O(n1241));
  orx  g1143(.A(n2331), .B(n227), .O(n1242));
  orx  g1144(.A(pi27), .B(n199), .O(n1243));
  orx  g1145(.A(pi27), .B(n214), .O(n1244));
  orx  g1146(.A(n2524), .B(n2360), .O(n1245));
  orx  g1147(.A(pi28), .B(n704), .O(n1246));
  orx  g1148(.A(n2421), .B(n705), .O(n1247));
  orx  g1149(.A(n709), .B(n710), .O(n1248));
  orx  g1150(.A(n713), .B(n714), .O(n1249));
  orx  g1151(.A(n715), .B(n716), .O(n1250));
  orx  g1152(.A(n717), .B(n718), .O(n1251));
  orx  g1153(.A(n719), .B(n720), .O(n1252));
  orx  g1154(.A(n721), .B(n722), .O(n1253));
  orx  g1155(.A(n2331), .B(n2531), .O(n1254));
  orx  g1156(.A(pi27), .B(n283), .O(n1255));
  orx  g1157(.A(pi28), .B(n280), .O(n1256));
  orx  g1158(.A(n2421), .B(n725), .O(n1257));
  orx  g1159(.A(n729), .B(n730), .O(n1258));
  orx  g1160(.A(n731), .B(n732), .O(n1259));
  orx  g1161(.A(n2331), .B(n2455), .O(n1260));
  orx  g1162(.A(pi28), .B(n733), .O(n1261));
  orx  g1163(.A(pi28), .B(n221), .O(n1262));
  orx  g1164(.A(n2422), .B(n289), .O(n1263));
  orx  g1165(.A(n738), .B(n739), .O(n1264));
  orx  g1166(.A(n2331), .B(n198), .O(n1265));
  orx  g1167(.A(pi27), .B(n288), .O(n1266));
  orx  g1168(.A(n2329), .B(n2532), .O(n1267));
  orx  g1169(.A(pi27), .B(n287), .O(n1268));
  orx  g1170(.A(pi28), .B(n741), .O(n1269));
  orx  g1171(.A(n2422), .B(n742), .O(n1270));
  orx  g1172(.A(n746), .B(n747), .O(n1271));
  orx  g1173(.A(n748), .B(n749), .O(n1272));
  orx  g1174(.A(n750), .B(n751), .O(n1273));
  orx  g1175(.A(n752), .B(n753), .O(n1274));
  orx  g1176(.A(n754), .B(n755), .O(n1275));
  orx  g1177(.A(n756), .B(n757), .O(n1276));
  orx  g1178(.A(n758), .B(n759), .O(n1277));
  orx  g1179(.A(n760), .B(n761), .O(n1278));
  orx  g1180(.A(pi27), .B(n237), .O(n1279));
  orx  g1181(.A(n2330), .B(n2531), .O(n1280));
  orx  g1182(.A(pi28), .B(n193), .O(n1281));
  orx  g1183(.A(n2422), .B(n762), .O(n1282));
  orx  g1184(.A(n766), .B(n767), .O(n1283));
  orx  g1185(.A(n770), .B(n771), .O(n1284));
  orx  g1186(.A(n772), .B(n773), .O(n1285));
  orx  g1187(.A(n776), .B(n777), .O(n1286));
  orx  g1188(.A(n778), .B(n779), .O(n1287));
  orx  g1189(.A(n780), .B(n781), .O(n1288));
  orx  g1190(.A(n782), .B(n783), .O(n1289));
  orx  g1191(.A(n784), .B(n785), .O(n1290));
  orx  g1192(.A(pi27), .B(n2307), .O(n1291));
  orx  g1193(.A(n2522), .B(n2359), .O(n1292));
  orx  g1194(.A(n2374), .B(n2344), .O(n1293));
  orx  g1195(.A(pi27), .B(n2589), .O(n1294));
  orx  g1196(.A(pi28), .B(n786), .O(n1295));
  orx  g1197(.A(n2422), .B(n787), .O(n1296));
  orx  g1198(.A(n791), .B(n792), .O(n1297));
  orx  g1199(.A(n2376), .B(n2312), .O(n1298));
  orx  g1200(.A(pi30), .B(n2317), .O(n1299));
  orx  g1201(.A(n794), .B(n795), .O(n1300));
  orx  g1202(.A(n796), .B(n797), .O(n1301));
  orx  g1203(.A(n800), .B(n801), .O(n1302));
  orx  g1204(.A(n804), .B(n805), .O(n1303));
  orx  g1205(.A(n806), .B(n807), .O(n1304));
  orx  g1206(.A(n808), .B(n809), .O(n1305));
  orx  g1207(.A(n2328), .B(n2454), .O(n1306));
  orx  g1208(.A(pi28), .B(n2498), .O(n1307));
  orx  g1209(.A(n2330), .B(n230), .O(n1308));
  orx  g1210(.A(pi27), .B(n2520), .O(n1309));
  orx  g1211(.A(pi28), .B(n811), .O(n1310));
  orx  g1212(.A(n2423), .B(n300), .O(n1311));
  orx  g1213(.A(n815), .B(n816), .O(n1312));
  orx  g1214(.A(n817), .B(n818), .O(n1313));
  orx  g1215(.A(n819), .B(n820), .O(n1314));
  orx  g1216(.A(n821), .B(n822), .O(n1315));
  orx  g1217(.A(n823), .B(n824), .O(n1316));
  orx  g1218(.A(n825), .B(n826), .O(n1317));
  orx  g1219(.A(n827), .B(n828), .O(n1318));
  orx  g1220(.A(n829), .B(n830), .O(n1319));
  orx  g1221(.A(n2319), .B(n2405), .O(n1320));
  orx  g1222(.A(pi30), .B(n2274), .O(n1321));
  orx  g1223(.A(n2329), .B(n2543), .O(n1322));
  orx  g1224(.A(pi27), .B(n831), .O(n1323));
  orx  g1225(.A(n2523), .B(n2360), .O(n1324));
  orx  g1226(.A(pi27), .B(n2578), .O(n1325));
  orx  g1227(.A(pi28), .B(n832), .O(n1326));
  orx  g1228(.A(n2423), .B(n833), .O(n1327));
  orx  g1229(.A(n2423), .B(n193), .O(n1328));
  orx  g1230(.A(pi28), .B(n218), .O(n1329));
  orx  g1231(.A(n840), .B(n841), .O(n1330));
  orx  g1232(.A(n842), .B(n843), .O(n1331));
  orx  g1233(.A(n844), .B(n845), .O(n1332));
  orx  g1234(.A(n846), .B(n847), .O(n1333));
  orx  g1235(.A(pi27), .B(pi29), .O(n1334));
  orx  g1236(.A(n2327), .B(n2516), .O(n1335));
  orx  g1237(.A(pi30), .B(n2277), .O(n1336));
  orx  g1238(.A(n2373), .B(n2312), .O(n1337));
  orx  g1239(.A(n2329), .B(n2532), .O(n1338));
  orx  g1240(.A(pi27), .B(n849), .O(n1339));
  orx  g1241(.A(pi28), .B(n848), .O(n1340));
  orx  g1242(.A(n2423), .B(n850), .O(n1341));
  orx  g1243(.A(n854), .B(n855), .O(n1342));
  orx  g1244(.A(n856), .B(n857), .O(n1343));
  orx  g1245(.A(n858), .B(n859), .O(n1344));
  orx  g1246(.A(n860), .B(n861), .O(n1345));
  orx  g1247(.A(n862), .B(n863), .O(n1346));
  orx  g1248(.A(n864), .B(n865), .O(n1347));
  orx  g1249(.A(pi27), .B(n234), .O(n1348));
  orx  g1250(.A(n2587), .B(n2360), .O(n1349));
  orx  g1251(.A(pi27), .B(n233), .O(n1350));
  orx  g1252(.A(n2524), .B(n2360), .O(n1351));
  orx  g1253(.A(pi28), .B(n866), .O(n1352));
  orx  g1254(.A(n2424), .B(n867), .O(n1353));
  orx  g1255(.A(n871), .B(n872), .O(n1354));
  orx  g1256(.A(n873), .B(n874), .O(n1355));
  orx  g1257(.A(n875), .B(n876), .O(n1356));
  orx  g1258(.A(n880), .B(n881), .O(n1357));
  orx  g1259(.A(n882), .B(n883), .O(n1358));
  orx  g1260(.A(n884), .B(n885), .O(n1359));
  orx  g1261(.A(pi28), .B(n264), .O(n1360));
  orx  g1262(.A(n2424), .B(n312), .O(n1361));
  orx  g1263(.A(n891), .B(n892), .O(n1362));
  orx  g1264(.A(n893), .B(n894), .O(n1363));
  orx  g1265(.A(n896), .B(n897), .O(n1364));
  orx  g1266(.A(n900), .B(n901), .O(n1365));
  orx  g1267(.A(n902), .B(n903), .O(n1366));
  orx  g1268(.A(n904), .B(n905), .O(n1367));
  orx  g1269(.A(pi28), .B(n906), .O(n1368));
  orx  g1270(.A(n2424), .B(n316), .O(n1369));
  orx  g1271(.A(n910), .B(n911), .O(n1370));
  orx  g1272(.A(n912), .B(n913), .O(n1371));
  orx  g1273(.A(n914), .B(n915), .O(n1372));
  orx  g1274(.A(n916), .B(n917), .O(n1373));
  orx  g1275(.A(n918), .B(n919), .O(n1374));
  orx  g1276(.A(n920), .B(n921), .O(n1375));
  orx  g1277(.A(n922), .B(n923), .O(n1376));
  orx  g1278(.A(pi27), .B(n2572), .O(n1377));
  orx  g1279(.A(n2327), .B(n201), .O(n1378));
  orx  g1280(.A(pi27), .B(n2520), .O(n1379));
  orx  g1281(.A(n2257), .B(n2346), .O(n1380));
  orx  g1282(.A(pi28), .B(n924), .O(n1381));
  orx  g1283(.A(n2424), .B(n925), .O(n1382));
  orx  g1284(.A(n929), .B(n930), .O(n1383));
  orx  g1285(.A(n931), .B(n932), .O(n1384));
  orx  g1286(.A(n933), .B(n934), .O(n1385));
  orx  g1287(.A(n935), .B(n936), .O(n1386));
  orx  g1288(.A(n937), .B(n938), .O(n1387));
  orx  g1289(.A(n2328), .B(n2586), .O(n1388));
  orx  g1290(.A(pi27), .B(n2551), .O(n1389));
  orx  g1291(.A(n2328), .B(n2532), .O(n1390));
  orx  g1292(.A(pi27), .B(n220), .O(n1391));
  orx  g1293(.A(pi28), .B(n939), .O(n1392));
  orx  g1294(.A(n2425), .B(n940), .O(n1393));
  orx  g1295(.A(n944), .B(n945), .O(n1394));
  orx  g1296(.A(n946), .B(n947), .O(n1395));
  orx  g1297(.A(n948), .B(n949), .O(n1396));
  orx  g1298(.A(n950), .B(n951), .O(n1397));
  orx  g1299(.A(n952), .B(n953), .O(n1398));
  orx  g1300(.A(n954), .B(n955), .O(n1399));
  orx  g1301(.A(n956), .B(n957), .O(n1400));
  orx  g1302(.A(pi27), .B(n215), .O(n1401));
  orx  g1303(.A(n2326), .B(n211), .O(n1402));
  orx  g1304(.A(pi28), .B(n958), .O(n1403));
  orx  g1305(.A(n2425), .B(n326), .O(n1404));
  orx  g1306(.A(n962), .B(n963), .O(n1405));
  orx  g1307(.A(n964), .B(n965), .O(n1406));
  orx  g1308(.A(n966), .B(n967), .O(n1407));
  orx  g1309(.A(n968), .B(n969), .O(n1408));
  orx  g1310(.A(n970), .B(n971), .O(n1409));
  orx  g1311(.A(n972), .B(n973), .O(n1410));
  orx  g1312(.A(n974), .B(n975), .O(n1411));
  orx  g1313(.A(pi28), .B(n229), .O(n1412));
  orx  g1314(.A(n2588), .B(n2453), .O(n1413));
  orx  g1315(.A(pi27), .B(n976), .O(n1414));
  orx  g1316(.A(n2328), .B(n329), .O(n1415));
  orx  g1317(.A(n980), .B(n981), .O(n1416));
  orx  g1318(.A(n982), .B(n983), .O(n1417));
  orx  g1319(.A(n985), .B(n984), .O(n1418));
  orx  g1320(.A(n987), .B(n986), .O(n1419));
  orx  g1321(.A(n988), .B(n989), .O(n1420));
  orx  g1322(.A(n990), .B(n991), .O(n1421));
  orx  g1323(.A(n2589), .B(n2361), .O(n1422));
  orx  g1324(.A(pi27), .B(n2552), .O(n1423));
  orx  g1325(.A(pi27), .B(n2603), .O(n1424));
  orx  g1326(.A(n2327), .B(n2562), .O(n1425));
  orx  g1327(.A(pi28), .B(n992), .O(n1426));
  orx  g1328(.A(n2425), .B(n993), .O(n1427));
  orx  g1329(.A(n998), .B(n997), .O(n1428));
  orx  g1330(.A(n1000), .B(n999), .O(n1429));
  orx  g1331(.A(n1001), .B(n1002), .O(n1430));
  orx  g1332(.A(n1004), .B(n1003), .O(n1431));
  orx  g1333(.A(n1005), .B(n1006), .O(n1432));
  orx  g1334(.A(n1007), .B(n1008), .O(n1433));
  orx  g1335(.A(n1009), .B(n1010), .O(n1434));
  orx  g1336(.A(pi27), .B(n2275), .O(n1435));
  orx  g1337(.A(n2326), .B(n283), .O(n1436));
  orx  g1338(.A(n2425), .B(n1165), .O(n1437));
  orx  g1339(.A(pi28), .B(n1011), .O(n1438));
  orx  g1340(.A(pi27), .B(n2320), .O(n1439));
  orx  g1341(.A(n2511), .B(n2306), .O(n1440));
  andx g1342(.A(n1972), .B(pi30), .O(n1441));
  orx  g1343(.A(n2264), .B(n2297), .O(n1442));
  orx  g1344(.A(n2612), .B(n2591), .O(n1443));
  orx  g1345(.A(n2268), .B(pi29), .O(n1444));
  andx g1346(.A(n1444), .B(pi25), .O(n1445));
  orx  g1347(.A(n2609), .B(n2306), .O(n1446));
  andx g1348(.A(n2306), .B(pi29), .O(n1447));
  andx g1349(.A(n1486), .B(pi30), .O(n1448));
  andx g1350(.A(n1936), .B(n2444), .O(n1449));
  orx  g1351(.A(n2591), .B(pi29), .O(n1450));
  andx g1352(.A(n1559), .B(n1964), .O(n1451));
  andx g1353(.A(n1992), .B(n1991), .O(n1452));
  andx g1354(.A(n2600), .B(n2389), .O(n1453));
  andx g1355(.A(n1993), .B(n2484), .O(n1454));
  orx  g1356(.A(n1454), .B(n2262), .O(n1455));
  andx g1357(.A(n1994), .B(n2484), .O(n1456));
  orx  g1358(.A(n1456), .B(n2295), .O(n1457));
  orx  g1359(.A(n2327), .B(n2318), .O(n1458));
  orx  g1360(.A(pi31), .B(n2335), .O(n1459));
  orx  g1361(.A(pi31), .B(pi27), .O(n1460));
  orx  g1362(.A(n2591), .B(n2297), .O(n1461));
  orx  g1363(.A(n2271), .B(n2671), .O(n1462));
  orx  g1364(.A(n2293), .B(n2270), .O(n1463));
  orx  g1365(.A(n2267), .B(n2604), .O(n1464));
  andx g1366(.A(n2497), .B(n2225), .O(n1465));
  orx  g1367(.A(pi29), .B(n2272), .O(n1466));
  orx  g1368(.A(n2271), .B(n2604), .O(n1467));
  orx  g1369(.A(pi31), .B(pi29), .O(n1468));
  orx  g1370(.A(n2263), .B(n2604), .O(n1469));
  andx g1371(.A(n2260), .B(n1988), .O(n1470));
  orx  g1372(.A(n2376), .B(n2592), .O(n1471));
  orx  g1373(.A(n2377), .B(n1462), .O(n1472));
  andx g1374(.A(n2402), .B(n2484), .O(n1473));
  orx  g1375(.A(n1571), .B(n1572), .O(n1474));
  orx  g1376(.A(n1561), .B(n1562), .O(n1475));
  orx  g1377(.A(n348), .B(n1598), .O(n1476));
  orx  g1378(.A(n1795), .B(n1878), .O(n1477));
  orx  g1379(.A(n1788), .B(n1565), .O(n1478));
  orx  g1380(.A(n1837), .B(n1899), .O(n1479));
  orx  g1381(.A(n1917), .B(n798), .O(n1480));
  orx  g1382(.A(n2301), .B(n2671), .O(n1481));
  andx g1383(.A(n1587), .B(n1971), .O(n1482));
  orx  g1384(.A(n1565), .B(n1566), .O(n1483));
  andx g1385(.A(n1588), .B(n2485), .O(n1484));
  orx  g1386(.A(n1590), .B(n1589), .O(n1485));
  orx  g1387(.A(n1612), .B(n1613), .O(n1486));
  orx  g1388(.A(n1603), .B(n1899), .O(n1487));
  orx  g1389(.A(n1599), .B(n1600), .O(n1488));
  orx  g1390(.A(n1591), .B(n1595), .O(n1489));
  andx g1391(.A(n1615), .B(n2485), .O(n1490));
  orx  g1392(.A(n1617), .B(n1616), .O(n1491));
  andx g1393(.A(n1633), .B(n2389), .O(n1492));
  orx  g1394(.A(n1625), .B(n1645), .O(n1493));
  orx  g1395(.A(n1623), .B(n1624), .O(n1494));
  andx g1396(.A(n1481), .B(n2300), .O(n1495));
  andx g1397(.A(n1974), .B(n2389), .O(n1496));
  andx g1398(.A(n1634), .B(n2485), .O(n1497));
  orx  g1399(.A(n1636), .B(n1635), .O(n1498));
  orx  g1400(.A(n1671), .B(n1658), .O(n1499));
  orx  g1401(.A(n1649), .B(n1573), .O(n1500));
  orx  g1402(.A(n1899), .B(n1648), .O(n1501));
  orx  g1403(.A(n1644), .B(n1645), .O(n1502));
  andx g1404(.A(pi29), .B(n2320), .O(n1503));
  andx g1405(.A(n1661), .B(n1657), .O(n1504));
  orx  g1406(.A(n1663), .B(n1662), .O(n1505));
  orx  g1407(.A(n1742), .B(n1683), .O(n1506));
  andx g1408(.A(n2621), .B(n1977), .O(n1507));
  andx g1409(.A(n1685), .B(n2485), .O(n1508));
  orx  g1410(.A(n1687), .B(n1686), .O(n1509));
  andx g1411(.A(n1704), .B(n2389), .O(n1510));
  orx  g1412(.A(n1695), .B(n1624), .O(n1511));
  andx g1413(.A(n1705), .B(n2486), .O(n1512));
  orx  g1414(.A(n1707), .B(n1706), .O(n1513));
  orx  g1415(.A(n1742), .B(n1726), .O(n1514));
  andx g1416(.A(n1728), .B(n2486), .O(n1515));
  orx  g1417(.A(n1730), .B(n1729), .O(n1516));
  orx  g1418(.A(n1742), .B(n1743), .O(n1517));
  andx g1419(.A(pi31), .B(n2486), .O(n1518));
  andx g1420(.A(n1557), .B(n1745), .O(n1519));
  orx  g1421(.A(n1747), .B(n1746), .O(n1520));
  andx g1422(.A(n1966), .B(n1083), .O(n1521));
  andx g1423(.A(n1765), .B(n2486), .O(n1522));
  orx  g1424(.A(n1767), .B(n1766), .O(n1523));
  andx g1425(.A(n1783), .B(n2487), .O(n1524));
  orx  g1426(.A(n1785), .B(n1784), .O(n1525));
  andx g1427(.A(n1807), .B(n2487), .O(n1526));
  orx  g1428(.A(n1809), .B(n1808), .O(n1527));
  andx g1429(.A(pi29), .B(pi31), .O(n1528));
  andx g1430(.A(n1980), .B(n1468), .O(n1529));
  andx g1431(.A(n1828), .B(n2487), .O(n1530));
  orx  g1432(.A(n1830), .B(n1829), .O(n1531));
  andx g1433(.A(n1834), .B(n2553), .O(n1532));
  andx g1434(.A(n1849), .B(n2487), .O(n1533));
  orx  g1435(.A(n1851), .B(n1850), .O(n1534));
  andx g1436(.A(n2601), .B(n2390), .O(n1535));
  andx g1437(.A(n1869), .B(n2488), .O(n1536));
  orx  g1438(.A(n1871), .B(n1870), .O(n1537));
  andx g1439(.A(n1981), .B(n2304), .O(n1538));
  andx g1440(.A(n1887), .B(n2488), .O(n1539));
  orx  g1441(.A(n1889), .B(n1888), .O(n1540));
  andx g1442(.A(n1983), .B(n1463), .O(n1541));
  andx g1443(.A(n2508), .B(n1982), .O(n1542));
  orx  g1444(.A(n1612), .B(n1890), .O(n1543));
  andx g1445(.A(n1906), .B(n2488), .O(n1544));
  orx  g1446(.A(n1908), .B(n1907), .O(n1545));
  andx g1447(.A(n1927), .B(n2488), .O(n1546));
  orx  g1448(.A(n1929), .B(n1928), .O(n1547));
  andx g1449(.A(n1987), .B(n1986), .O(n1548));
  andx g1450(.A(n1941), .B(n1939), .O(n1549));
  orx  g1451(.A(n1942), .B(n1943), .O(n1550));
  andx g1452(.A(n1558), .B(n1951), .O(n1551));
  orx  g1453(.A(n1955), .B(n1954), .O(n1552));
  andx g1454(.A(n1961), .B(n1960), .O(n1553));
  orx  g1455(.A(n1963), .B(n1962), .O(n1554));
  orx  g1456(.A(n2591), .B(n2292), .O(n1555));
  orx  g1457(.A(n2306), .B(n2297), .O(n1556));
  andx g1458(.A(n1968), .B(n2489), .O(n1557));
  andx g1459(.A(n1953), .B(n2489), .O(n1558));
  andx g1460(.A(pi28), .B(n2489), .O(n1559));
  orx  g1461(.A(n2426), .B(n2497), .O(n1560));
  andx g1462(.A(pi29), .B(n2270), .O(n1561));
  andx g1463(.A(n2591), .B(n2671), .O(n1562));
  andx g1464(.A(pi30), .B(pi27), .O(n1563));
  andx g1465(.A(n1475), .B(n2390), .O(n1564));
  andx g1466(.A(n2299), .B(n2292), .O(n1565));
  andx g1467(.A(n2590), .B(pi29), .O(n1566));
  andx g1468(.A(n1483), .B(n2390), .O(n1567));
  andx g1469(.A(n2518), .B(pi30), .O(n1568));
  andx g1470(.A(n1995), .B(n2445), .O(n1569));
  andx g1471(.A(n1996), .B(pi28), .O(n1570));
  andx g1472(.A(pi31), .B(n2355), .O(n1571));
  andx g1473(.A(pi27), .B(n2318), .O(n1572));
  andx g1474(.A(n1458), .B(n2293), .O(n1573));
  andx g1475(.A(n2301), .B(pi29), .O(n1574));
  orx  g1476(.A(pi29), .B(n2264), .O(n1575));
  andx g1477(.A(n1998), .B(n2391), .O(n1576));
  andx g1478(.A(n2597), .B(pi30), .O(n1577));
  orx  g1479(.A(pi29), .B(n2673), .O(n1578));
  andx g1480(.A(n1970), .B(n2391), .O(n1579));
  andx g1481(.A(n2596), .B(pi30), .O(n1580));
  andx g1482(.A(n1999), .B(n2444), .O(n1581));
  andx g1483(.A(n2000), .B(pi28), .O(n1582));
  andx g1484(.A(n1997), .B(n2469), .O(n1583));
  andx g1485(.A(n2001), .B(pi25), .O(n1584));
  andx g1486(.A(n2004), .B(n2003), .O(n1585));
  andx g1487(.A(n2006), .B(n2005), .O(n1586));
  andx g1488(.A(n2008), .B(n2007), .O(n1587));
  andx g1489(.A(n2010), .B(n2009), .O(n1588));
  andx g1490(.A(n2002), .B(n2295), .O(n1589));
  andx g1491(.A(n1484), .B(pi26), .O(n1590));
  andx g1492(.A(n2291), .B(n2318), .O(n1591));
  andx g1493(.A(pi29), .B(n2263), .O(n1592));
  andx g1494(.A(n1440), .B(n2391), .O(n1593));
  andx g1495(.A(n2011), .B(pi30), .O(n1594));
  andx g1496(.A(n2301), .B(pi29), .O(n1595));
  andx g1497(.A(n2012), .B(n2444), .O(n1596));
  andx g1498(.A(n1973), .B(pi28), .O(n1597));
  andx g1499(.A(pi29), .B(n2318), .O(n1598));
  andx g1500(.A(pi29), .B(pi31), .O(n1599));
  andx g1501(.A(n2305), .B(n2266), .O(n1600));
  andx g1502(.A(n1476), .B(n2391), .O(n1601));
  andx g1503(.A(n1488), .B(pi30), .O(n1602));
  andx g1504(.A(pi29), .B(n2319), .O(n1603));
  andx g1505(.A(n1487), .B(n2392), .O(n1604));
  andx g1506(.A(n1442), .B(pi30), .O(n1605));
  andx g1507(.A(n2014), .B(n2445), .O(n1606));
  andx g1508(.A(n2015), .B(pi28), .O(n1607));
  andx g1509(.A(n2013), .B(n2489), .O(n1608));
  andx g1510(.A(n2016), .B(pi25), .O(n1609));
  andx g1511(.A(n2019), .B(n2018), .O(n1610));
  andx g1512(.A(n2021), .B(n2020), .O(n1611));
  andx g1513(.A(n2265), .B(n2356), .O(n1612));
  andx g1514(.A(pi29), .B(n2272), .O(n1613));
  andx g1515(.A(n2023), .B(n2022), .O(n1614));
  andx g1516(.A(n2025), .B(n2024), .O(n1615));
  andx g1517(.A(n2017), .B(n2286), .O(n1616));
  andx g1518(.A(n1490), .B(pi26), .O(n1617));
  andx g1519(.A(n2306), .B(pi29), .O(n1618));
  andx g1520(.A(n2026), .B(n2392), .O(n1619));
  andx g1521(.A(n1495), .B(pi30), .O(n1620));
  andx g1522(.A(n2027), .B(n2447), .O(n1621));
  andx g1523(.A(n1496), .B(pi28), .O(n1622));
  andx g1524(.A(pi29), .B(n2354), .O(n1623));
  andx g1525(.A(n2301), .B(n2293), .O(n1624));
  andx g1526(.A(pi29), .B(pi31), .O(n1625));
  andx g1527(.A(n1481), .B(n2392), .O(n1626));
  andx g1528(.A(n1493), .B(pi30), .O(n1627));
  andx g1529(.A(n1975), .B(n2444), .O(n1628));
  andx g1530(.A(n2029), .B(pi28), .O(n1629));
  andx g1531(.A(n2028), .B(n2486), .O(n1630));
  andx g1532(.A(n2030), .B(pi25), .O(n1631));
  andx g1533(.A(n2033), .B(n2032), .O(n1632));
  andx g1534(.A(n2035), .B(n2034), .O(n1633));
  andx g1535(.A(n2037), .B(n2036), .O(n1634));
  andx g1536(.A(n2031), .B(n2287), .O(n1635));
  andx g1537(.A(n1497), .B(pi26), .O(n1636));
  andx g1538(.A(pi29), .B(n2264), .O(n1637));
  andx g1539(.A(n1503), .B(n2466), .O(n1638));
  andx g1540(.A(n2038), .B(pi25), .O(n1639));
  andx g1541(.A(n2506), .B(pi25), .O(n1640));
  andx g1542(.A(n1976), .B(n2484), .O(n1641));
  andx g1543(.A(n2039), .B(n2393), .O(n1642));
  andx g1544(.A(n2040), .B(pi30), .O(n1643));
  andx g1545(.A(n2267), .B(pi29), .O(n1644));
  andx g1546(.A(n2264), .B(n2265), .O(n1645));
  andx g1547(.A(n2607), .B(n2651), .O(n1646));
  andx g1548(.A(n1502), .B(pi25), .O(n1647));
  andx g1549(.A(n2305), .B(pi29), .O(n1648));
  andx g1550(.A(pi29), .B(pi31), .O(n1649));
  andx g1551(.A(n1501), .B(n2492), .O(n1650));
  andx g1552(.A(n1500), .B(pi25), .O(n1651));
  andx g1553(.A(n2042), .B(n2393), .O(n1652));
  andx g1554(.A(n2043), .B(pi30), .O(n1653));
  andx g1555(.A(n2041), .B(n2448), .O(n1654));
  andx g1556(.A(n2044), .B(pi28), .O(n1655));
  orx  g1557(.A(pi30), .B(n2455), .O(n1656));
  andx g1558(.A(n2047), .B(n2046), .O(n1657));
  andx g1559(.A(n2305), .B(pi29), .O(n1658));
  andx g1560(.A(n2049), .B(n2048), .O(n1659));
  andx g1561(.A(n2051), .B(n2050), .O(n1660));
  andx g1562(.A(n2053), .B(n2052), .O(n1661));
  andx g1563(.A(n2045), .B(n2295), .O(n1662));
  andx g1564(.A(n1504), .B(pi26), .O(n1663));
  andx g1565(.A(n2297), .B(n2394), .O(n1664));
  andx g1566(.A(n1443), .B(pi30), .O(n1665));
  andx g1567(.A(n2507), .B(pi30), .O(n1666));
  andx g1568(.A(n2620), .B(n2394), .O(n1667));
  andx g1569(.A(n2054), .B(n2448), .O(n1668));
  andx g1570(.A(n2055), .B(pi28), .O(n1669));
  andx g1571(.A(pi29), .B(n2356), .O(n1670));
  andx g1572(.A(n2272), .B(n2671), .O(n1671));
  andx g1573(.A(n2519), .B(n2393), .O(n1672));
  andx g1574(.A(n2057), .B(pi30), .O(n1673));
  andx g1575(.A(pi29), .B(n2300), .O(n1674));
  andx g1576(.A(n2590), .B(n2265), .O(n1675));
  andx g1577(.A(n1474), .B(pi29), .O(n1676));
  andx g1578(.A(n2059), .B(n2395), .O(n1677));
  andx g1579(.A(n2060), .B(pi30), .O(n1678));
  andx g1580(.A(n2058), .B(n2445), .O(n1679));
  andx g1581(.A(n2061), .B(pi28), .O(n1680));
  andx g1582(.A(n2056), .B(n2483), .O(n1681));
  andx g1583(.A(n2062), .B(pi25), .O(n1682));
  andx g1584(.A(n2591), .B(pi29), .O(n1683));
  andx g1585(.A(n2065), .B(n2064), .O(n1684));
  andx g1586(.A(n2067), .B(n2066), .O(n1685));
  andx g1587(.A(n2063), .B(n2633), .O(n1686));
  andx g1588(.A(n1508), .B(pi26), .O(n1687));
  andx g1589(.A(n1476), .B(pi30), .O(n1688));
  andx g1590(.A(n2514), .B(n2395), .O(n1689));
  andx g1591(.A(pi29), .B(n1458), .O(n1690));
  andx g1592(.A(pi30), .B(n1083), .O(n1691));
  andx g1593(.A(n2069), .B(n2393), .O(n1692));
  andx g1594(.A(n2068), .B(n2443), .O(n1693));
  andx g1595(.A(n2070), .B(pi28), .O(n1694));
  andx g1596(.A(pi29), .B(pi27), .O(n1695));
  andx g1597(.A(pi30), .B(n2512), .O(n1696));
  andx g1598(.A(n1499), .B(n2395), .O(n1697));
  andx g1599(.A(n1978), .B(n2446), .O(n1698));
  andx g1600(.A(n2072), .B(pi28), .O(n1699));
  andx g1601(.A(n2071), .B(n2490), .O(n1700));
  andx g1602(.A(n2073), .B(pi25), .O(n1701));
  andx g1603(.A(n2076), .B(n2075), .O(n1702));
  andx g1604(.A(n2078), .B(n2077), .O(n1703));
  andx g1605(.A(n2079), .B(n1462), .O(n1704));
  andx g1606(.A(n2081), .B(n2080), .O(n1705));
  andx g1607(.A(n2074), .B(n2285), .O(n1706));
  andx g1608(.A(n1512), .B(pi26), .O(n1707));
  andx g1609(.A(pi31), .B(n2396), .O(n1708));
  andx g1610(.A(n2301), .B(pi30), .O(n1709));
  andx g1611(.A(pi29), .B(n2272), .O(n1710));
  andx g1612(.A(pi29), .B(n2394), .O(n1711));
  andx g1613(.A(n2083), .B(pi30), .O(n1712));
  andx g1614(.A(n2082), .B(n2449), .O(n1713));
  andx g1615(.A(n2084), .B(pi28), .O(n1714));
  andx g1616(.A(n1489), .B(pi30), .O(n1715));
  andx g1617(.A(n2304), .B(n2396), .O(n1716));
  andx g1618(.A(n2299), .B(pi29), .O(n1717));
  andx g1619(.A(n1483), .B(pi30), .O(n1718));
  andx g1620(.A(n2087), .B(n2396), .O(n1719));
  andx g1621(.A(n2086), .B(n2447), .O(n1720));
  andx g1622(.A(n2088), .B(pi28), .O(n1721));
  andx g1623(.A(n2085), .B(n2484), .O(n1722));
  andx g1624(.A(n2089), .B(pi25), .O(n1723));
  orx  g1625(.A(n2609), .B(n2267), .O(n1724));
  andx g1626(.A(n2092), .B(n2091), .O(n1725));
  andx g1627(.A(pi29), .B(n1459), .O(n1726));
  andx g1628(.A(n2094), .B(n2093), .O(n1727));
  andx g1629(.A(n2096), .B(n2095), .O(n1728));
  andx g1630(.A(n2090), .B(n2284), .O(n1729));
  andx g1631(.A(n1515), .B(pi26), .O(n1730));
  andx g1632(.A(n1518), .B(n2392), .O(n1731));
  andx g1633(.A(n1979), .B(pi30), .O(n1732));
  andx g1634(.A(n2591), .B(pi29), .O(n1733));
  andx g1635(.A(n1464), .B(n2490), .O(n1734));
  andx g1636(.A(n2098), .B(pi25), .O(n1735));
  andx g1637(.A(n2508), .B(n2490), .O(n1736));
  andx g1638(.A(n2617), .B(pi25), .O(n1737));
  andx g1639(.A(n2099), .B(n2397), .O(n1738));
  andx g1640(.A(n2100), .B(pi30), .O(n1739));
  andx g1641(.A(n2097), .B(n2450), .O(n1740));
  andx g1642(.A(n2101), .B(pi28), .O(n1741));
  andx g1643(.A(pi27), .B(n2291), .O(n1742));
  andx g1644(.A(pi29), .B(n2270), .O(n1743));
  andx g1645(.A(n2104), .B(n2103), .O(n1744));
  andx g1646(.A(n2106), .B(n2105), .O(n1745));
  andx g1647(.A(n2102), .B(n2284), .O(n1746));
  andx g1648(.A(n1519), .B(pi26), .O(n1747));
  andx g1649(.A(pi25), .B(n2319), .O(n1748));
  andx g1650(.A(n2306), .B(n2491), .O(n1749));
  orx  g1651(.A(pi29), .B(n2299), .O(n1750));
  andx g1652(.A(n2597), .B(pi25), .O(n1751));
  andx g1653(.A(n2595), .B(n2490), .O(n1752));
  andx g1654(.A(n2107), .B(n2397), .O(n1753));
  andx g1655(.A(n2108), .B(pi30), .O(n1754));
  andx g1656(.A(n2622), .B(pi25), .O(n1755));
  andx g1657(.A(n1517), .B(n2491), .O(n1756));
  andx g1658(.A(n2267), .B(n2491), .O(n1757));
  andx g1659(.A(n1521), .B(pi25), .O(n1758));
  andx g1660(.A(n2110), .B(n2395), .O(n1759));
  andx g1661(.A(n2111), .B(pi30), .O(n1760));
  andx g1662(.A(n2109), .B(n2446), .O(n1761));
  andx g1663(.A(n2112), .B(pi28), .O(n1762));
  andx g1664(.A(n2115), .B(n2114), .O(n1763));
  andx g1665(.A(n2117), .B(n2116), .O(n1764));
  andx g1666(.A(n2119), .B(n2118), .O(n1765));
  andx g1667(.A(n2113), .B(n2261), .O(n1766));
  andx g1668(.A(n1522), .B(pi26), .O(n1767));
  andx g1669(.A(n2623), .B(n2450), .O(n1768));
  andx g1670(.A(pi28), .B(n2614), .O(n1769));
  andx g1671(.A(n2610), .B(n2447), .O(n1770));
  andx g1672(.A(n2605), .B(pi28), .O(n1771));
  andx g1673(.A(n2120), .B(n2398), .O(n1772));
  andx g1674(.A(n2121), .B(pi30), .O(n1773));
  andx g1675(.A(pi28), .B(n1461), .O(n1774));
  andx g1676(.A(n2007), .B(n2451), .O(n1775));
  andx g1677(.A(n1969), .B(n2396), .O(n1776));
  andx g1678(.A(n2123), .B(pi30), .O(n1777));
  andx g1679(.A(n2122), .B(n2492), .O(n1778));
  andx g1680(.A(n2124), .B(pi25), .O(n1779));
  orx  g1681(.A(n1459), .B(pi29), .O(n1780));
  andx g1682(.A(n2127), .B(n2126), .O(n1781));
  andx g1683(.A(n2129), .B(n2128), .O(n1782));
  andx g1684(.A(n2131), .B(n2130), .O(n1783));
  andx g1685(.A(n2125), .B(n2287), .O(n1784));
  andx g1686(.A(n1524), .B(pi26), .O(n1785));
  andx g1687(.A(pi25), .B(n1460), .O(n1786));
  andx g1688(.A(n2087), .B(n2491), .O(n1787));
  andx g1689(.A(pi29), .B(n2272), .O(n1788));
  andx g1690(.A(n2511), .B(n2492), .O(n1789));
  andx g1691(.A(n2616), .B(pi25), .O(n1790));
  andx g1692(.A(n2132), .B(n2398), .O(n1791));
  andx g1693(.A(n2133), .B(pi30), .O(n1792));
  andx g1694(.A(pi31), .B(n2492), .O(n1793));
  andx g1695(.A(pi25), .B(n2263), .O(n1794));
  andx g1696(.A(pi29), .B(n2493), .O(n1795));
  andx g1697(.A(n2553), .B(n2590), .O(n1796));
  andx g1698(.A(n1477), .B(n2135), .O(n1797));
  andx g1699(.A(n2297), .B(n2492), .O(n1798));
  andx g1700(.A(n1500), .B(pi25), .O(n1799));
  andx g1701(.A(n2136), .B(n2397), .O(n1800));
  andx g1702(.A(n2137), .B(pi30), .O(n1801));
  andx g1703(.A(n2134), .B(n2447), .O(n1802));
  andx g1704(.A(n2138), .B(pi28), .O(n1803));
  andx g1705(.A(n2141), .B(n2140), .O(n1804));
  andx g1706(.A(n2143), .B(n2142), .O(n1805));
  andx g1707(.A(n2145), .B(n2144), .O(n1806));
  andx g1708(.A(n2147), .B(n2146), .O(n1807));
  andx g1709(.A(n2139), .B(n2262), .O(n1808));
  andx g1710(.A(n1526), .B(pi26), .O(n1809));
  andx g1711(.A(n2299), .B(pi29), .O(n1810));
  andx g1712(.A(n2148), .B(n2493), .O(n1811));
  andx g1713(.A(n1528), .B(pi25), .O(n1812));
  andx g1714(.A(n2149), .B(n2399), .O(n1813));
  andx g1715(.A(n1529), .B(pi30), .O(n1814));
  andx g1716(.A(n2007), .B(n2151), .O(n1815));
  andx g1717(.A(n2268), .B(n2493), .O(n1816));
  andx g1718(.A(n1815), .B(pi25), .O(n1817));
  andx g1719(.A(pi25), .B(pi27), .O(n1818));
  andx g1720(.A(n2299), .B(n2494), .O(n1819));
  andx g1721(.A(n1477), .B(pi31), .O(n1820));
  andx g1722(.A(n2153), .B(n2553), .O(n1821));
  andx g1723(.A(n2152), .B(n2399), .O(n1822));
  andx g1724(.A(n2154), .B(pi30), .O(n1823));
  andx g1725(.A(n2150), .B(n2445), .O(n1824));
  andx g1726(.A(n2155), .B(pi28), .O(n1825));
  andx g1727(.A(n2158), .B(n2157), .O(n1826));
  andx g1728(.A(n2160), .B(n2159), .O(n1827));
  andx g1729(.A(n2162), .B(n2161), .O(n1828));
  andx g1730(.A(n2156), .B(n2294), .O(n1829));
  andx g1731(.A(n1530), .B(pi26), .O(n1830));
  andx g1732(.A(pi29), .B(pi27), .O(n1831));
  andx g1733(.A(n2606), .B(n2493), .O(n1832));
  andx g1734(.A(n2163), .B(pi25), .O(n1833));
  andx g1735(.A(n2166), .B(n2165), .O(n1834));
  andx g1736(.A(n2164), .B(n2399), .O(n1835));
  andx g1737(.A(n1532), .B(pi30), .O(n1836));
  andx g1738(.A(n2301), .B(pi29), .O(n1837));
  andx g1739(.A(n1469), .B(n2494), .O(n1838));
  andx g1740(.A(n1479), .B(pi25), .O(n1839));
  andx g1741(.A(n1474), .B(pi29), .O(n1840));
  andx g1742(.A(n2596), .B(pi25), .O(n1841));
  andx g1743(.A(n2169), .B(n2494), .O(n1842));
  andx g1744(.A(n2168), .B(n2397), .O(n1843));
  andx g1745(.A(n2170), .B(pi30), .O(n1844));
  andx g1746(.A(n2167), .B(n2448), .O(n1845));
  andx g1747(.A(n2171), .B(pi28), .O(n1846));
  andx g1748(.A(n2174), .B(n2173), .O(n1847));
  andx g1749(.A(n2176), .B(n2175), .O(n1848));
  andx g1750(.A(n2178), .B(n2177), .O(n1849));
  andx g1751(.A(n2172), .B(n2260), .O(n1850));
  andx g1752(.A(n1533), .B(pi26), .O(n1851));
  andx g1753(.A(n2506), .B(pi30), .O(n1852));
  andx g1754(.A(n2057), .B(n2400), .O(n1853));
  andx g1755(.A(pi29), .B(pi27), .O(n1854));
  andx g1756(.A(n1478), .B(pi30), .O(n1855));
  andx g1757(.A(n2180), .B(n2400), .O(n1856));
  andx g1758(.A(n2179), .B(n2451), .O(n1857));
  andx g1759(.A(n2181), .B(pi28), .O(n1858));
  andx g1760(.A(pi29), .B(n2319), .O(n1859));
  andx g1761(.A(n2509), .B(pi30), .O(n1860));
  andx g1762(.A(n2183), .B(n2394), .O(n1861));
  andx g1763(.A(pi30), .B(n2266), .O(n1862));
  andx g1764(.A(n2517), .B(n2400), .O(n1863));
  andx g1765(.A(n2184), .B(n2448), .O(n1864));
  andx g1766(.A(n2185), .B(pi28), .O(n1865));
  andx g1767(.A(n2182), .B(n2495), .O(n1866));
  andx g1768(.A(n2186), .B(pi25), .O(n1867));
  andx g1769(.A(n2189), .B(n2188), .O(n1868));
  andx g1770(.A(n2191), .B(n2190), .O(n1869));
  andx g1771(.A(n2187), .B(n2286), .O(n1870));
  andx g1772(.A(n1536), .B(pi26), .O(n1871));
  andx g1773(.A(n1443), .B(n2494), .O(n1872));
  andx g1774(.A(n1506), .B(pi25), .O(n1873));
  andx g1775(.A(n1538), .B(n2398), .O(n1874));
  andx g1776(.A(n2192), .B(pi30), .O(n1875));
  andx g1777(.A(n1488), .B(n2495), .O(n1876));
  andx g1778(.A(n1486), .B(pi25), .O(n1877));
  andx g1779(.A(pi25), .B(n2291), .O(n1878));
  andx g1780(.A(n2059), .B(n2495), .O(n1879));
  andx g1781(.A(n2194), .B(n2400), .O(n1880));
  andx g1782(.A(n2195), .B(pi30), .O(n1881));
  andx g1783(.A(n2193), .B(n2446), .O(n1882));
  andx g1784(.A(n2196), .B(pi28), .O(n1883));
  andx g1785(.A(n2199), .B(n2198), .O(n1884));
  orx  g1786(.A(n2590), .B(pi29), .O(n1885));
  andx g1787(.A(n2201), .B(n2200), .O(n1886));
  andx g1788(.A(n2203), .B(n2202), .O(n1887));
  andx g1789(.A(n2197), .B(n2260), .O(n1888));
  andx g1790(.A(n1539), .B(pi26), .O(n1889));
  andx g1791(.A(n2268), .B(pi29), .O(n1890));
  andx g1792(.A(n2304), .B(n2449), .O(n1891));
  andx g1793(.A(n1543), .B(pi28), .O(n1892));
  andx g1794(.A(n2510), .B(n2451), .O(n1893));
  andx g1795(.A(n2060), .B(pi28), .O(n1894));
  andx g1796(.A(n2204), .B(n2401), .O(n1895));
  andx g1797(.A(n2205), .B(pi30), .O(n1896));
  andx g1798(.A(pi28), .B(n2321), .O(n1897));
  andx g1799(.A(n2300), .B(n2449), .O(n1898));
  andx g1800(.A(n1474), .B(n2265), .O(n1899));
  andx g1801(.A(n2207), .B(pi29), .O(n1900));
  andx g1802(.A(n2208), .B(n2398), .O(n1901));
  andx g1803(.A(n1542), .B(pi30), .O(n1902));
  andx g1804(.A(n2206), .B(n2496), .O(n1903));
  andx g1805(.A(n2209), .B(pi25), .O(n1904));
  andx g1806(.A(n2212), .B(n2211), .O(n1905));
  andx g1807(.A(n2214), .B(n2213), .O(n1906));
  andx g1808(.A(n2210), .B(n2259), .O(n1907));
  andx g1809(.A(n1544), .B(pi26), .O(n1908));
  andx g1810(.A(pi30), .B(n1463), .O(n1909));
  andx g1811(.A(n2304), .B(n2401), .O(n1910));
  andx g1812(.A(n2215), .B(n2451), .O(n1911));
  andx g1813(.A(n1984), .B(pi28), .O(n1912));
  andx g1814(.A(n2615), .B(pi30), .O(n1913));
  andx g1815(.A(n1985), .B(n2401), .O(n1914));
  andx g1816(.A(pi30), .B(pi31), .O(n1915));
  andx g1817(.A(n2271), .B(n2399), .O(n1916));
  andx g1818(.A(pi29), .B(n2401), .O(n1917));
  andx g1819(.A(n1480), .B(n2356), .O(n1918));
  andx g1820(.A(n2218), .B(n2534), .O(n1919));
  andx g1821(.A(n2217), .B(n2449), .O(n1920));
  andx g1822(.A(n2219), .B(pi28), .O(n1921));
  andx g1823(.A(n2216), .B(n2495), .O(n1922));
  andx g1824(.A(n2220), .B(pi25), .O(n1923));
  andx g1825(.A(n2223), .B(n2222), .O(n1924));
  andx g1826(.A(n2225), .B(n2224), .O(n1925));
  andx g1827(.A(n2226), .B(n2145), .O(n1926));
  andx g1828(.A(n2228), .B(n2227), .O(n1927));
  andx g1829(.A(n2221), .B(n2295), .O(n1928));
  andx g1830(.A(n1546), .B(pi26), .O(n1929));
  andx g1831(.A(pi28), .B(n1462), .O(n1930));
  andx g1832(.A(n2304), .B(n2446), .O(n1931));
  andx g1833(.A(pi28), .B(n1464), .O(n1932));
  andx g1834(.A(n2619), .B(n2450), .O(n1933));
  andx g1835(.A(n2229), .B(n2633), .O(n1934));
  andx g1836(.A(n2230), .B(pi26), .O(n1935));
  andx g1837(.A(n2232), .B(n2233), .O(n1936));
  andx g1838(.A(n2231), .B(n2402), .O(n1937));
  andx g1839(.A(n1548), .B(pi30), .O(n1938));
  andx g1840(.A(n2236), .B(n2235), .O(n1939));
  andx g1841(.A(n2238), .B(n2237), .O(n1940));
  andx g1842(.A(n2240), .B(n2239), .O(n1941));
  andx g1843(.A(n2234), .B(n2496), .O(n1942));
  andx g1844(.A(n1549), .B(pi25), .O(n1943));
  andx g1845(.A(n1989), .B(n2452), .O(n1944));
  andx g1846(.A(pi28), .B(n1472), .O(n1945));
  andx g1847(.A(n2515), .B(pi30), .O(n1946));
  andx g1848(.A(n2536), .B(n2450), .O(n1947));
  andx g1849(.A(n2242), .B(pi28), .O(n1948));
  andx g1850(.A(n2241), .B(n2496), .O(n1949));
  andx g1851(.A(n2243), .B(pi25), .O(n1950));
  andx g1852(.A(n2246), .B(n2245), .O(n1951));
  orx  g1853(.A(n2608), .B(n2406), .O(n1952));
  andx g1854(.A(n2248), .B(n2247), .O(n1953));
  andx g1855(.A(n2244), .B(n2262), .O(n1954));
  andx g1856(.A(n1551), .B(pi26), .O(n1955));
  andx g1857(.A(n1989), .B(n2496), .O(n1956));
  andx g1858(.A(pi25), .B(n1471), .O(n1957));
  andx g1859(.A(n2249), .B(n2452), .O(n1958));
  andx g1860(.A(n1990), .B(pi28), .O(n1959));
  andx g1861(.A(n2252), .B(n2251), .O(n1960));
  andx g1862(.A(n2254), .B(n2253), .O(n1961));
  andx g1863(.A(n2250), .B(n2262), .O(n1962));
  andx g1864(.A(n1553), .B(pi26), .O(n1963));
  andx g1865(.A(n2256), .B(n2255), .O(n1964));
  orx  g1866(.A(pi29), .B(n2305), .O(n1965));
  orx  g1867(.A(n2265), .B(n2268), .O(n1966));
  orx  g1868(.A(n2291), .B(n2263), .O(n1967));
  orx  g1869(.A(n2374), .B(n2433), .O(n1968));
  orx  g1870(.A(n2427), .B(n1468), .O(n1969));
  orx  g1871(.A(n2511), .B(n2268), .O(n1970));
  orx  g1872(.A(n2594), .B(n2406), .O(n1971));
  orx  g1873(.A(pi29), .B(n2321), .O(n1972));
  orx  g1874(.A(n1489), .B(n1441), .O(n1973));
  orx  g1875(.A(n1458), .B(pi29), .O(n1974));
  orx  g1876(.A(n1494), .B(pi30), .O(n1975));
  orx  g1877(.A(pi29), .B(pi27), .O(n1976));
  orx  g1878(.A(n2599), .B(n2406), .O(n1977));
  orx  g1879(.A(n1511), .B(n2406), .O(n1978));
  orx  g1880(.A(n1446), .B(n1445), .O(n1979));
  orx  g1881(.A(n1447), .B(n2497), .O(n1980));
  orx  g1882(.A(n1502), .B(n2497), .O(n1981));
  orx  g1883(.A(n2598), .B(n2453), .O(n1982));
  orx  g1884(.A(n2592), .B(n2455), .O(n1983));
  orx  g1885(.A(n1448), .B(n2297), .O(n1984));
  orx  g1886(.A(n2511), .B(n2299), .O(n1985));
  orx  g1887(.A(n1449), .B(n2286), .O(n1986));
  orx  g1888(.A(n2515), .B(n2668), .O(n1987));
  orx  g1889(.A(n2513), .B(n2453), .O(n1988));
  orx  g1890(.A(n2304), .B(pi30), .O(n1989));
  orx  g1891(.A(n2535), .B(n2498), .O(n1990));
  orx  g1892(.A(n1451), .B(n2294), .O(n1991));
  orx  g1893(.A(n1472), .B(n1560), .O(n1992));
  orx  g1894(.A(n1453), .B(n2455), .O(n1993));
  orx  g1895(.A(n1471), .B(n2453), .O(n1994));
  orx  g1896(.A(n1563), .B(n1564), .O(n1995));
  orx  g1897(.A(n1567), .B(n1568), .O(n1996));
  orx  g1898(.A(n1569), .B(n1570), .O(n1997));
  orx  g1899(.A(n1573), .B(n1574), .O(n1998));
  orx  g1900(.A(n1576), .B(n1577), .O(n1999));
  orx  g1901(.A(n1579), .B(n1580), .O(n2000));
  orx  g1902(.A(n1581), .B(n1582), .O(n2001));
  orx  g1903(.A(n1583), .B(n1584), .O(n2002));
  orx  g1904(.A(pi29), .B(n2300), .O(n2003));
  orx  g1905(.A(n2305), .B(n2266), .O(n2004));
  orx  g1906(.A(pi30), .B(n1481), .O(n2005));
  orx  g1907(.A(n2376), .B(n1585), .O(n2006));
  orx  g1908(.A(pi27), .B(n2292), .O(n2007));
  orx  g1909(.A(pi29), .B(n2264), .O(n2008));
  orx  g1910(.A(pi28), .B(n1586), .O(n2009));
  orx  g1911(.A(n2430), .B(n1482), .O(n2010));
  orx  g1912(.A(n1591), .B(n1592), .O(n2011));
  orx  g1913(.A(n1593), .B(n1594), .O(n2012));
  orx  g1914(.A(n1596), .B(n1597), .O(n2013));
  orx  g1915(.A(n1601), .B(n1602), .O(n2014));
  orx  g1916(.A(n1604), .B(n1605), .O(n2015));
  orx  g1917(.A(n1606), .B(n1607), .O(n2016));
  orx  g1918(.A(n1608), .B(n1609), .O(n2017));
  orx  g1919(.A(n2326), .B(n2293), .O(n2018));
  orx  g1920(.A(pi29), .B(n2270), .O(n2019));
  orx  g1921(.A(pi30), .B(n2514), .O(n2020));
  orx  g1922(.A(n2375), .B(n1610), .O(n2021));
  orx  g1923(.A(n2594), .B(n2406), .O(n2022));
  orx  g1924(.A(pi30), .B(n1486), .O(n2023));
  orx  g1925(.A(pi28), .B(n1611), .O(n2024));
  orx  g1926(.A(n2427), .B(n1614), .O(n2025));
  orx  g1927(.A(n1562), .B(n1618), .O(n2026));
  orx  g1928(.A(n1619), .B(n1620), .O(n2027));
  orx  g1929(.A(n1621), .B(n1622), .O(n2028));
  orx  g1930(.A(n1626), .B(n1627), .O(n2029));
  orx  g1931(.A(n1628), .B(n1629), .O(n2030));
  orx  g1932(.A(n1630), .B(n1631), .O(n2031));
  orx  g1933(.A(n2375), .B(n2512), .O(n2032));
  orx  g1934(.A(pi30), .B(n2517), .O(n2033));
  orx  g1935(.A(pi27), .B(pi29), .O(n2034));
  orx  g1936(.A(n2266), .B(n1460), .O(n2035));
  orx  g1937(.A(pi28), .B(n1632), .O(n2036));
  orx  g1938(.A(n2430), .B(n1492), .O(n2037));
  orx  g1939(.A(n1742), .B(n1637), .O(n2038));
  orx  g1940(.A(n1638), .B(n1639), .O(n2039));
  orx  g1941(.A(n1640), .B(n1641), .O(n2040));
  orx  g1942(.A(n1642), .B(n1643), .O(n2041));
  orx  g1943(.A(n1646), .B(n1647), .O(n2042));
  orx  g1944(.A(n1650), .B(n1651), .O(n2043));
  orx  g1945(.A(n1652), .B(n1653), .O(n2044));
  orx  g1946(.A(n1654), .B(n1655), .O(n2045));
  orx  g1947(.A(n2533), .B(n2498), .O(n2046));
  orx  g1948(.A(n1465), .B(n1656), .O(n2047));
  orx  g1949(.A(n2305), .B(n2407), .O(n2048));
  orx  g1950(.A(pi30), .B(n1499), .O(n2049));
  orx  g1951(.A(pi30), .B(n2270), .O(n2050));
  orx  g1952(.A(n2373), .B(n2592), .O(n2051));
  orx  g1953(.A(pi28), .B(n1659), .O(n2052));
  orx  g1954(.A(n2428), .B(n1660), .O(n2053));
  orx  g1955(.A(n1664), .B(n1665), .O(n2054));
  orx  g1956(.A(n1666), .B(n1667), .O(n2055));
  orx  g1957(.A(n1668), .B(n1669), .O(n2056));
  orx  g1958(.A(n1670), .B(n1671), .O(n2057));
  orx  g1959(.A(n1672), .B(n1673), .O(n2058));
  orx  g1960(.A(n1674), .B(n1675), .O(n2059));
  orx  g1961(.A(n1742), .B(n1676), .O(n2060));
  orx  g1962(.A(n1677), .B(n1678), .O(n2061));
  orx  g1963(.A(n1679), .B(n1680), .O(n2062));
  orx  g1964(.A(n1681), .B(n1682), .O(n2063));
  orx  g1965(.A(n2375), .B(n2509), .O(n2064));
  orx  g1966(.A(pi30), .B(n1506), .O(n2065));
  orx  g1967(.A(pi28), .B(n1684), .O(n2066));
  orx  g1968(.A(n2430), .B(n1507), .O(n2067));
  orx  g1969(.A(n1688), .B(n1689), .O(n2068));
  orx  g1970(.A(n1690), .B(n1624), .O(n2069));
  orx  g1971(.A(n1691), .B(n1692), .O(n2070));
  orx  g1972(.A(n1693), .B(n1694), .O(n2071));
  orx  g1973(.A(n1696), .B(n1697), .O(n2072));
  orx  g1974(.A(n1698), .B(n1699), .O(n2073));
  orx  g1975(.A(n1700), .B(n1701), .O(n2074));
  orx  g1976(.A(pi31), .B(n2266), .O(n2075));
  orx  g1977(.A(pi29), .B(n2300), .O(n2076));
  orx  g1978(.A(pi30), .B(n2606), .O(n2077));
  orx  g1979(.A(n2375), .B(n1702), .O(n2078));
  orx  g1980(.A(pi29), .B(n2590), .O(n2079));
  orx  g1981(.A(pi28), .B(n1703), .O(n2080));
  orx  g1982(.A(n2426), .B(n1510), .O(n2081));
  orx  g1983(.A(n1708), .B(n1709), .O(n2082));
  orx  g1984(.A(n1573), .B(n1710), .O(n2083));
  orx  g1985(.A(n1711), .B(n1712), .O(n2084));
  orx  g1986(.A(n1713), .B(n1714), .O(n2085));
  orx  g1987(.A(n1715), .B(n1716), .O(n2086));
  orx  g1988(.A(n348), .B(n1717), .O(n2087));
  orx  g1989(.A(n1718), .B(n1719), .O(n2088));
  orx  g1990(.A(n1720), .B(n1721), .O(n2089));
  orx  g1991(.A(n1722), .B(n1723), .O(n2090));
  orx  g1992(.A(pi30), .B(n2598), .O(n2091));
  orx  g1993(.A(n2373), .B(n1724), .O(n2092));
  orx  g1994(.A(n2599), .B(n2408), .O(n2093));
  orx  g1995(.A(pi30), .B(n1514), .O(n2094));
  orx  g1996(.A(pi28), .B(n1725), .O(n2095));
  orx  g1997(.A(n2426), .B(n1727), .O(n2096));
  orx  g1998(.A(n1731), .B(n1732), .O(n2097));
  orx  g1999(.A(n1591), .B(n1733), .O(n2098));
  orx  g2000(.A(n1734), .B(n1735), .O(n2099));
  orx  g2001(.A(n1736), .B(n1737), .O(n2100));
  orx  g2002(.A(n1738), .B(n1739), .O(n2101));
  orx  g2003(.A(n1740), .B(n1741), .O(n2102));
  orx  g2004(.A(n2374), .B(n1483), .O(n2103));
  orx  g2005(.A(pi30), .B(n1517), .O(n2104));
  orx  g2006(.A(n1461), .B(n2454), .O(n2105));
  orx  g2007(.A(pi28), .B(n1744), .O(n2106));
  orx  g2008(.A(n1748), .B(n1749), .O(n2107));
  orx  g2009(.A(n1751), .B(n1752), .O(n2108));
  orx  g2010(.A(n1753), .B(n1754), .O(n2109));
  orx  g2011(.A(n1755), .B(n1756), .O(n2110));
  orx  g2012(.A(n1757), .B(n1758), .O(n2111));
  orx  g2013(.A(n1759), .B(n1760), .O(n2112));
  orx  g2014(.A(n1761), .B(n1762), .O(n2113));
  orx  g2015(.A(pi30), .B(n1517), .O(n2114));
  orx  g2016(.A(n2608), .B(n2407), .O(n2115));
  orx  g2017(.A(pi30), .B(n2297), .O(n2116));
  orx  g2018(.A(n2594), .B(n2407), .O(n2117));
  orx  g2019(.A(pi28), .B(n1763), .O(n2118));
  orx  g2020(.A(n2428), .B(n1764), .O(n2119));
  orx  g2021(.A(n1768), .B(n1769), .O(n2120));
  orx  g2022(.A(n1770), .B(n1771), .O(n2121));
  orx  g2023(.A(n1772), .B(n1773), .O(n2122));
  orx  g2024(.A(n1774), .B(n1775), .O(n2123));
  orx  g2025(.A(n1776), .B(n1777), .O(n2124));
  orx  g2026(.A(n1778), .B(n1779), .O(n2125));
  orx  g2027(.A(pi28), .B(n2618), .O(n2126));
  orx  g2028(.A(n2430), .B(n1780), .O(n2127));
  orx  g2029(.A(pi28), .B(n2361), .O(n2128));
  orx  g2030(.A(n2431), .B(n2592), .O(n2129));
  orx  g2031(.A(pi30), .B(n1781), .O(n2130));
  orx  g2032(.A(n2374), .B(n1782), .O(n2131));
  orx  g2033(.A(n1786), .B(n1787), .O(n2132));
  orx  g2034(.A(n1789), .B(n1790), .O(n2133));
  orx  g2035(.A(n1791), .B(n1792), .O(n2134));
  orx  g2036(.A(n1793), .B(n1794), .O(n2135));
  orx  g2037(.A(n1796), .B(n1797), .O(n2136));
  orx  g2038(.A(n1798), .B(n1799), .O(n2137));
  orx  g2039(.A(n1800), .B(n1801), .O(n2138));
  orx  g2040(.A(n1802), .B(n1803), .O(n2139));
  orx  g2041(.A(pi31), .B(pi30), .O(n2140));
  orx  g2042(.A(n2305), .B(n2407), .O(n2141));
  orx  g2043(.A(pi29), .B(n2270), .O(n2142));
  orx  g2044(.A(n2292), .B(n1804), .O(n2143));
  orx  g2045(.A(pi30), .B(n2263), .O(n2144));
  orx  g2046(.A(n2373), .B(n2592), .O(n2145));
  orx  g2047(.A(pi28), .B(n1805), .O(n2146));
  orx  g2048(.A(n2428), .B(n1806), .O(n2147));
  orx  g2049(.A(n1810), .B(n1899), .O(n2148));
  orx  g2050(.A(n1811), .B(n1812), .O(n2149));
  orx  g2051(.A(n1813), .B(n1814), .O(n2150));
  orx  g2052(.A(pi29), .B(n2361), .O(n2151));
  orx  g2053(.A(n1816), .B(n1817), .O(n2152));
  orx  g2054(.A(n1818), .B(n1819), .O(n2153));
  orx  g2055(.A(n1820), .B(n1821), .O(n2154));
  orx  g2056(.A(n1822), .B(n1823), .O(n2155));
  orx  g2057(.A(n1824), .B(n1825), .O(n2156));
  orx  g2058(.A(pi30), .B(n2361), .O(n2157));
  orx  g2059(.A(n2515), .B(n2407), .O(n2158));
  orx  g2060(.A(n2372), .B(n2592), .O(n2159));
  orx  g2061(.A(pi30), .B(n1478), .O(n2160));
  orx  g2062(.A(pi28), .B(n1826), .O(n2161));
  orx  g2063(.A(n2426), .B(n1827), .O(n2162));
  orx  g2064(.A(n1831), .B(n348), .O(n2163));
  orx  g2065(.A(n1832), .B(n1833), .O(n2164));
  orx  g2066(.A(pi25), .B(n2361), .O(n2165));
  orx  g2067(.A(pi27), .B(n2498), .O(n2166));
  orx  g2068(.A(n1835), .B(n1836), .O(n2167));
  orx  g2069(.A(n1838), .B(n1839), .O(n2168));
  orx  g2070(.A(n1565), .B(n1840), .O(n2169));
  orx  g2071(.A(n1841), .B(n1842), .O(n2170));
  orx  g2072(.A(n1843), .B(n1844), .O(n2171));
  orx  g2073(.A(n1845), .B(n1846), .O(n2172));
  orx  g2074(.A(n2371), .B(n1476), .O(n2173));
  orx  g2075(.A(pi30), .B(n2612), .O(n2174));
  orx  g2076(.A(n2372), .B(n2592), .O(n2175));
  orx  g2077(.A(pi30), .B(n2605), .O(n2176));
  orx  g2078(.A(pi28), .B(n1847), .O(n2177));
  orx  g2079(.A(n2429), .B(n1848), .O(n2178));
  orx  g2080(.A(n1852), .B(n1853), .O(n2179));
  orx  g2081(.A(n1854), .B(n1675), .O(n2180));
  orx  g2082(.A(n1855), .B(n1856), .O(n2181));
  orx  g2083(.A(n1857), .B(n1858), .O(n2182));
  orx  g2084(.A(n1859), .B(n1624), .O(n2183));
  orx  g2085(.A(n1860), .B(n1861), .O(n2184));
  orx  g2086(.A(n1862), .B(n1863), .O(n2185));
  orx  g2087(.A(n1864), .B(n1865), .O(n2186));
  orx  g2088(.A(n1866), .B(n1867), .O(n2187));
  orx  g2089(.A(pi30), .B(n2511), .O(n2188));
  orx  g2090(.A(n2371), .B(n1479), .O(n2189));
  orx  g2091(.A(pi28), .B(n1868), .O(n2190));
  orx  g2092(.A(n2431), .B(n1535), .O(n2191));
  orx  g2093(.A(n1872), .B(n1873), .O(n2192));
  orx  g2094(.A(n1874), .B(n1875), .O(n2193));
  orx  g2095(.A(n1876), .B(n1877), .O(n2194));
  orx  g2096(.A(n1878), .B(n1879), .O(n2195));
  orx  g2097(.A(n1880), .B(n1881), .O(n2196));
  orx  g2098(.A(n1882), .B(n1883), .O(n2197));
  orx  g2099(.A(pi29), .B(pi30), .O(n2198));
  orx  g2100(.A(n2372), .B(n1467), .O(n2199));
  orx  g2101(.A(n2372), .B(n2592), .O(n2200));
  orx  g2102(.A(pi30), .B(n1885), .O(n2201));
  orx  g2103(.A(pi28), .B(n1884), .O(n2202));
  orx  g2104(.A(n2427), .B(n1886), .O(n2203));
  orx  g2105(.A(n1891), .B(n1892), .O(n2204));
  orx  g2106(.A(n1893), .B(n1894), .O(n2205));
  orx  g2107(.A(n1895), .B(n1896), .O(n2206));
  orx  g2108(.A(n1897), .B(n1898), .O(n2207));
  orx  g2109(.A(n1899), .B(n1900), .O(n2208));
  orx  g2110(.A(n1901), .B(n1902), .O(n2209));
  orx  g2111(.A(n1903), .B(n1904), .O(n2210));
  orx  g2112(.A(pi29), .B(pi28), .O(n2211));
  orx  g2113(.A(n1446), .B(n2453), .O(n2212));
  orx  g2114(.A(pi30), .B(n1905), .O(n2213));
  orx  g2115(.A(n2371), .B(n1541), .O(n2214));
  orx  g2116(.A(n1909), .B(n1910), .O(n2215));
  orx  g2117(.A(n1911), .B(n1912), .O(n2216));
  orx  g2118(.A(n1913), .B(n1914), .O(n2217));
  orx  g2119(.A(n1915), .B(n1916), .O(n2218));
  orx  g2120(.A(n1918), .B(n1919), .O(n2219));
  orx  g2121(.A(n1920), .B(n1921), .O(n2220));
  orx  g2122(.A(n1922), .B(n1923), .O(n2221));
  orx  g2123(.A(pi30), .B(n1476), .O(n2222));
  orx  g2124(.A(n2598), .B(n2408), .O(n2223));
  orx  g2125(.A(pi27), .B(pi29), .O(n2224));
  orx  g2126(.A(n2306), .B(n2293), .O(n2225));
  orx  g2127(.A(pi30), .B(n1925), .O(n2226));
  orx  g2128(.A(pi28), .B(n1924), .O(n2227));
  orx  g2129(.A(n2429), .B(n1926), .O(n2228));
  orx  g2130(.A(n1930), .B(n1931), .O(n2229));
  orx  g2131(.A(n1932), .B(n1933), .O(n2230));
  orx  g2132(.A(n1935), .B(n1934), .O(n2231));
  orx  g2133(.A(n2321), .B(n2265), .O(n2232));
  orx  g2134(.A(pi29), .B(n2356), .O(n2233));
  orx  g2135(.A(n1937), .B(n1938), .O(n2234));
  orx  g2136(.A(pi30), .B(n2260), .O(n2235));
  orx  g2137(.A(n2381), .B(n1470), .O(n2236));
  orx  g2138(.A(pi28), .B(n2266), .O(n2237));
  orx  g2139(.A(pi29), .B(n2454), .O(n2238));
  orx  g2140(.A(n2403), .B(n1517), .O(n2239));
  orx  g2141(.A(pi30), .B(n1940), .O(n2240));
  orx  g2142(.A(n1944), .B(n1945), .O(n2241));
  orx  g2143(.A(n625), .B(n1946), .O(n2242));
  orx  g2144(.A(n1947), .B(n1948), .O(n2243));
  orx  g2145(.A(n1949), .B(n1950), .O(n2244));
  orx  g2146(.A(n2427), .B(n2611), .O(n2245));
  orx  g2147(.A(pi28), .B(n1750), .O(n2246));
  orx  g2148(.A(n2669), .B(n2452), .O(n2247));
  orx  g2149(.A(pi28), .B(n1952), .O(n2248));
  orx  g2150(.A(n1956), .B(n1957), .O(n2249));
  orx  g2151(.A(n1958), .B(n1959), .O(n2250));
  orx  g2152(.A(pi28), .B(n2498), .O(n2251));
  orx  g2153(.A(n2429), .B(n1473), .O(n2252));
  orx  g2154(.A(n1443), .B(n2454), .O(n2253));
  orx  g2155(.A(pi28), .B(n2534), .O(n2254));
  orx  g2156(.A(n2599), .B(n2408), .O(n2255));
  orx  g2157(.A(pi30), .B(n1450), .O(n2256));
  invx g2158(.A(n1336), .O(n2257));
  invx g2159(.A(n2257), .O(n2258));
  invx g2160(.A(pi26), .O(n2259));
  invx g2161(.A(pi26), .O(n2260));
  invx g2162(.A(pi26), .O(n2261));
  invx g2163(.A(pi26), .O(n2262));
  invx g2164(.A(n1439), .O(n2263));
  invx g2165(.A(n1439), .O(n2264));
  invx g2166(.A(pi29), .O(n2265));
  invx g2167(.A(pi29), .O(n2266));
  invx g2168(.A(n1474), .O(n2267));
  invx g2169(.A(n2267), .O(n2268));
  invx g2170(.A(n1458), .O(n2269));
  invx g2171(.A(n2269), .O(n2270));
  invx g2172(.A(n1460), .O(n2271));
  invx g2173(.A(n2271), .O(n2272));
  invx g2174(.A(n190), .O(n2273));
  invx g2175(.A(n2273), .O(n2274));
  invx g2176(.A(n2273), .O(n2275));
  invx g2177(.A(n190), .O(n2276));
  invx g2178(.A(n190), .O(n2277));
  invx g2179(.A(n163), .O(n2278));
  invx g2180(.A(n2278), .O(n2279));
  invx g2181(.A(n2278), .O(n2280));
  invx g2182(.A(n2278), .O(n2281));
  invx g2183(.A(n2279), .O(n2282));
  invx g2184(.A(n163), .O(n2283));
  invx g2185(.A(pi26), .O(n2284));
  invx g2186(.A(pi26), .O(n2285));
  invx g2187(.A(pi26), .O(n2286));
  invx g2188(.A(pi26), .O(n2287));
  invx g2189(.A(n205), .O(n2288));
  invx g2190(.A(n2288), .O(n2289));
  invx g2191(.A(n2288), .O(n2290));
  invx g2192(.A(pi29), .O(n2291));
  invx g2193(.A(pi29), .O(n2292));
  invx g2194(.A(pi29), .O(n2293));
  invx g2195(.A(pi26), .O(n2294));
  invx g2196(.A(pi26), .O(n2295));
  bufx g2197(.A(n2298), .O(n2296));
  bufx g2198(.A(n2515), .O(n2297));
  bufx g2199(.A(n2726), .O(n2298));
  bufx g2200(.A(n2271), .O(n2299));
  bufx g2201(.A(n1459), .O(n2300));
  bufx g2202(.A(n2267), .O(n2301));
  bufx g2203(.A(n2602), .O(n2302));
  bufx g2204(.A(n2602), .O(n2303));
  bufx g2205(.A(n1466), .O(n2304));
  bufx g2206(.A(n1439), .O(n2305));
  bufx g2207(.A(n2590), .O(n2306));
  bufx g2208(.A(n2288), .O(n2307));
  bufx g2209(.A(n2288), .O(n2308));
  invx g2210(.A(n2322), .O(n2309));
  invx g2211(.A(n2322), .O(n2310));
  invx g2212(.A(n2322), .O(n2311));
  bufx g2213(.A(n2316), .O(n2312));
  bufx g2214(.A(n2316), .O(n2313));
  bufx g2215(.A(n164), .O(n2314));
  bufx g2216(.A(n164), .O(n2315));
  invx g2217(.A(n166), .O(n2316));
  invx g2218(.A(n2316), .O(n2317));
  invx g2219(.A(pi31), .O(n2318));
  invx g2220(.A(pi31), .O(n2319));
  invx g2221(.A(pi31), .O(n2320));
  invx g2222(.A(pi31), .O(n2321));
  invx g2223(.A(n2726), .O(n2322));
  invx g2224(.A(n2322), .O(n2323));
  invx g2225(.A(n2322), .O(n2324));
  invx g2226(.A(n2322), .O(n2325));
  invx g2227(.A(n2370), .O(n2326));
  invx g2228(.A(n2369), .O(n2327));
  invx g2229(.A(n2369), .O(n2328));
  invx g2230(.A(n2369), .O(n2329));
  invx g2231(.A(n2368), .O(n2330));
  invx g2232(.A(n2368), .O(n2331));
  invx g2233(.A(n2368), .O(n2332));
  invx g2234(.A(n2369), .O(n2333));
  invx g2235(.A(n2370), .O(n2334));
  invx g2236(.A(n2366), .O(n2335));
  invx g2237(.A(n2367), .O(n2336));
  invx g2238(.A(n2367), .O(n2337));
  invx g2239(.A(n2367), .O(n2338));
  invx g2240(.A(n2366), .O(n2339));
  invx g2241(.A(n2363), .O(n2340));
  invx g2242(.A(n2364), .O(n2341));
  invx g2243(.A(n2366), .O(n2342));
  invx g2244(.A(n2366), .O(n2343));
  invx g2245(.A(n2366), .O(n2344));
  invx g2246(.A(n2370), .O(n2345));
  invx g2247(.A(n2370), .O(n2346));
  invx g2248(.A(n2365), .O(n2347));
  invx g2249(.A(n2367), .O(n2348));
  invx g2250(.A(n2365), .O(n2349));
  invx g2251(.A(n2365), .O(n2350));
  invx g2252(.A(n2365), .O(n2351));
  invx g2253(.A(n2364), .O(n2352));
  invx g2254(.A(n2364), .O(n2353));
  invx g2255(.A(n2364), .O(n2354));
  invx g2256(.A(n2363), .O(n2355));
  invx g2257(.A(n2363), .O(n2356));
  invx g2258(.A(n2363), .O(n2357));
  invx g2259(.A(n2362), .O(n2358));
  invx g2260(.A(n2362), .O(n2359));
  invx g2261(.A(n2362), .O(n2360));
  invx g2262(.A(n2368), .O(n2361));
  invx g2263(.A(n2341), .O(n2362));
  invx g2264(.A(n2336), .O(n2363));
  invx g2265(.A(n2337), .O(n2364));
  invx g2266(.A(n2338), .O(n2365));
  invx g2267(.A(n2348), .O(n2366));
  invx g2268(.A(n2673), .O(n2367));
  invx g2269(.A(n2339), .O(n2368));
  invx g2270(.A(n2342), .O(n2369));
  invx g2271(.A(n2343), .O(n2370));
  invx g2272(.A(n2410), .O(n2371));
  invx g2273(.A(n2410), .O(n2372));
  invx g2274(.A(n2417), .O(n2373));
  invx g2275(.A(n2417), .O(n2374));
  invx g2276(.A(n2417), .O(n2375));
  invx g2277(.A(n2416), .O(n2376));
  invx g2278(.A(n2416), .O(n2377));
  invx g2279(.A(n2416), .O(n2378));
  invx g2280(.A(n2411), .O(n2379));
  invx g2281(.A(n2412), .O(n2380));
  invx g2282(.A(n2413), .O(n2381));
  invx g2283(.A(n2414), .O(n2382));
  invx g2284(.A(n2415), .O(n2383));
  invx g2285(.A(n2411), .O(n2384));
  invx g2286(.A(n2414), .O(n2385));
  invx g2287(.A(n2415), .O(n2386));
  invx g2288(.A(n2416), .O(n2387));
  invx g2289(.A(n2412), .O(n2388));
  invx g2290(.A(n2417), .O(n2389));
  invx g2291(.A(n2415), .O(n2390));
  invx g2292(.A(n2415), .O(n2391));
  invx g2293(.A(n2415), .O(n2392));
  invx g2294(.A(n2414), .O(n2393));
  invx g2295(.A(n2414), .O(n2394));
  invx g2296(.A(n2414), .O(n2395));
  invx g2297(.A(n2413), .O(n2396));
  invx g2298(.A(n2413), .O(n2397));
  invx g2299(.A(n2413), .O(n2398));
  invx g2300(.A(n2412), .O(n2399));
  invx g2301(.A(n2412), .O(n2400));
  invx g2302(.A(n2412), .O(n2401));
  invx g2303(.A(n2416), .O(n2402));
  invx g2304(.A(n2417), .O(n2403));
  invx g2305(.A(n2411), .O(n2404));
  invx g2306(.A(n2411), .O(n2405));
  invx g2307(.A(n2411), .O(n2406));
  invx g2308(.A(n2410), .O(n2407));
  invx g2309(.A(n2410), .O(n2408));
  invx g2310(.A(n2410), .O(n2409));
  invx g2311(.A(n2669), .O(n2410));
  invx g2312(.A(n2409), .O(n2411));
  invx g2313(.A(n2402), .O(n2412));
  invx g2314(.A(n2384), .O(n2413));
  invx g2315(.A(n2401), .O(n2414));
  invx g2316(.A(n2378), .O(n2415));
  invx g2317(.A(n2669), .O(n2416));
  invx g2318(.A(n2400), .O(n2417));
  invx g2319(.A(n2463), .O(n2418));
  invx g2320(.A(n2460), .O(n2419));
  invx g2321(.A(n2463), .O(n2420));
  invx g2322(.A(n2463), .O(n2421));
  invx g2323(.A(n2463), .O(n2422));
  invx g2324(.A(n2461), .O(n2423));
  invx g2325(.A(n2462), .O(n2424));
  invx g2326(.A(n2463), .O(n2425));
  invx g2327(.A(n2462), .O(n2426));
  invx g2328(.A(n2462), .O(n2427));
  invx g2329(.A(n2462), .O(n2428));
  invx g2330(.A(n2461), .O(n2429));
  invx g2331(.A(n2461), .O(n2430));
  invx g2332(.A(n2461), .O(n2431));
  invx g2333(.A(n2460), .O(n2432));
  invx g2334(.A(n2460), .O(n2433));
  invx g2335(.A(n2460), .O(n2434));
  invx g2336(.A(n2457), .O(n2435));
  invx g2337(.A(n2458), .O(n2436));
  invx g2338(.A(n2459), .O(n2437));
  invx g2339(.A(n2459), .O(n2438));
  invx g2340(.A(n2459), .O(n2439));
  invx g2341(.A(n2460), .O(n2440));
  invx g2342(.A(n2456), .O(n2441));
  invx g2343(.A(n2458), .O(n2442));
  invx g2344(.A(n2458), .O(n2443));
  invx g2345(.A(n2458), .O(n2444));
  invx g2346(.A(n2462), .O(n2445));
  invx g2347(.A(n2461), .O(n2446));
  invx g2348(.A(n2457), .O(n2447));
  invx g2349(.A(n2457), .O(n2448));
  invx g2350(.A(n2457), .O(n2449));
  invx g2351(.A(n2457), .O(n2450));
  invx g2352(.A(n2456), .O(n2451));
  invx g2353(.A(n2456), .O(n2452));
  invx g2354(.A(n2456), .O(n2453));
  invx g2355(.A(n2456), .O(n2454));
  invx g2356(.A(n2459), .O(n2455));
  invx g2357(.A(n2432), .O(n2456));
  invx g2358(.A(n2425), .O(n2457));
  invx g2359(.A(n2418), .O(n2458));
  invx g2360(.A(n2668), .O(n2459));
  invx g2361(.A(n2439), .O(n2460));
  invx g2362(.A(n2452), .O(n2461));
  invx g2363(.A(n2440), .O(n2462));
  invx g2364(.A(n2668), .O(n2463));
  invx g2365(.A(n2503), .O(n2464));
  invx g2366(.A(n2504), .O(n2465));
  invx g2367(.A(n2501), .O(n2466));
  invx g2368(.A(n2502), .O(n2467));
  invx g2369(.A(n2505), .O(n2468));
  invx g2370(.A(n2501), .O(n2469));
  invx g2371(.A(n2502), .O(n2470));
  invx g2372(.A(n2505), .O(n2471));
  invx g2373(.A(n2505), .O(n2472));
  invx g2374(.A(n2505), .O(n2473));
  invx g2375(.A(n2504), .O(n2474));
  invx g2376(.A(n2504), .O(n2475));
  invx g2377(.A(n2504), .O(n2476));
  invx g2378(.A(n2503), .O(n2477));
  invx g2379(.A(n2503), .O(n2478));
  invx g2380(.A(n2503), .O(n2479));
  invx g2381(.A(n2502), .O(n2480));
  invx g2382(.A(n2502), .O(n2481));
  invx g2383(.A(n2502), .O(n2482));
  invx g2384(.A(n2501), .O(n2483));
  invx g2385(.A(n2501), .O(n2484));
  invx g2386(.A(n2501), .O(n2485));
  invx g2387(.A(n2503), .O(n2486));
  invx g2388(.A(n2500), .O(n2487));
  invx g2389(.A(n2504), .O(n2488));
  invx g2390(.A(n2500), .O(n2489));
  invx g2391(.A(n2505), .O(n2490));
  invx g2392(.A(n2499), .O(n2491));
  invx g2393(.A(n2500), .O(n2492));
  invx g2394(.A(n2500), .O(n2493));
  invx g2395(.A(n2500), .O(n2494));
  invx g2396(.A(n2500), .O(n2495));
  invx g2397(.A(n2499), .O(n2496));
  invx g2398(.A(n2499), .O(n2497));
  invx g2399(.A(n2499), .O(n2498));
  invx g2400(.A(n2651), .O(n2499));
  invx g2401(.A(n2651), .O(n2500));
  invx g2402(.A(n2488), .O(n2501));
  invx g2403(.A(n2465), .O(n2502));
  invx g2404(.A(n2487), .O(n2503));
  invx g2405(.A(n2489), .O(n2504));
  invx g2406(.A(n2493), .O(n2505));
  invx g2407(.A(n1487), .O(n2506));
  invx g2408(.A(n1488), .O(n2507));
  invx g2409(.A(n1476), .O(n2508));
  invx g2410(.A(n1489), .O(n2509));
  invx g2411(.A(n1475), .O(n2510));
  invx g2412(.A(n1555), .O(n2511));
  invx g2413(.A(n1440), .O(n2512));
  invx g2414(.A(n1481), .O(n2513));
  invx g2415(.A(n1463), .O(n2514));
  invx g2416(.A(n1462), .O(n2515));
  invx g2417(.A(n170), .O(n2516));
  invx g2418(.A(n1556), .O(n2517));
  invx g2419(.A(n1461), .O(n2518));
  invx g2420(.A(n1442), .O(n2519));
  invx g2421(.A(n1015), .O(n2520));
  invx g2422(.A(n895), .O(n2521));
  invx g2423(.A(n338), .O(n2522));
  invx g2424(.A(n1146), .O(n2523));
  invx g2425(.A(n202), .O(n2524));
  invx g2426(.A(n199), .O(n2525));
  invx g2427(.A(n1018), .O(n2526));
  invx g2428(.A(n198), .O(n2527));
  invx g2429(.A(n196), .O(n2528));
  invx g2430(.A(n195), .O(n2529));
  invx g2431(.A(n194), .O(n2530));
  invx g2432(.A(n177), .O(n2531));
  invx g2433(.A(n167), .O(n2532));
  invx g2434(.A(n1656), .O(n2533));
  invx g2435(.A(n1480), .O(n2534));
  invx g2436(.A(n1472), .O(n2535));
  invx g2437(.A(n1471), .O(n2536));
  invx g2438(.A(n1031), .O(n2537));
  invx g2439(.A(n203), .O(n2538));
  invx g2440(.A(n1025), .O(n2539));
  invx g2441(.A(n546), .O(n2540));
  invx g2442(.A(n200), .O(n2541));
  invx g2443(.A(n171), .O(n2542));
  invx g2444(.A(n1024), .O(n2543));
  invx g2445(.A(n204), .O(n2544));
  invx g2446(.A(n173), .O(n2545));
  invx g2447(.A(n1019), .O(n2546));
  invx g2448(.A(n317), .O(n2547));
  invx g2449(.A(n318), .O(n2548));
  invx g2450(.A(n879), .O(n2549));
  invx g2451(.A(n313), .O(n2550));
  invx g2452(.A(n208), .O(n2551));
  invx g2453(.A(n301), .O(n2552));
  invx g2454(.A(n1477), .O(n2553));
  invx g2455(.A(n296), .O(n2554));
  invx g2456(.A(n297), .O(n2555));
  invx g2457(.A(n288), .O(n2556));
  invx g2458(.A(n283), .O(n2557));
  invx g2459(.A(n284), .O(n2558));
  invx g2460(.A(n697), .O(n2559));
  invx g2461(.A(n191), .O(n2560));
  invx g2462(.A(n169), .O(n2561));
  invx g2463(.A(n280), .O(n2562));
  invx g2464(.A(n277), .O(n2563));
  invx g2465(.A(n1212), .O(n2564));
  invx g2466(.A(n274), .O(n2565));
  invx g2467(.A(n261), .O(n2566));
  invx g2468(.A(n251), .O(n2567));
  invx g2469(.A(n253), .O(n2568));
  invx g2470(.A(n247), .O(n2569));
  invx g2471(.A(n242), .O(n2570));
  invx g2472(.A(n207), .O(n2571));
  invx g2473(.A(n243), .O(n2572));
  invx g2474(.A(n235), .O(n2573));
  invx g2475(.A(n237), .O(n2574));
  invx g2476(.A(n238), .O(n2575));
  invx g2477(.A(n236), .O(n2576));
  invx g2478(.A(n227), .O(n2577));
  invx g2479(.A(n228), .O(n2578));
  invx g2480(.A(n206), .O(n2579));
  invx g2481(.A(n219), .O(n2580));
  invx g2482(.A(n212), .O(n2581));
  invx g2483(.A(n213), .O(n2582));
  invx g2484(.A(n214), .O(n2583));
  invx g2485(.A(n215), .O(n2584));
  invx g2486(.A(n339), .O(n2585));
  invx g2487(.A(n336), .O(n2586));
  invx g2488(.A(n337), .O(n2587));
  invx g2489(.A(n201), .O(n2588));
  invx g2490(.A(n197), .O(n2589));
  invx g2491(.A(n1459), .O(n2590));
  invx g2492(.A(n2270), .O(n2591));
  invx g2493(.A(n1976), .O(n2592));
  invx g2494(.A(n193), .O(n2593));
  invx g2495(.A(n1965), .O(n2594));
  invx g2496(.A(n1750), .O(n2595));
  invx g2497(.A(n1578), .O(n2596));
  invx g2498(.A(n1575), .O(n2597));
  invx g2499(.A(n1468), .O(n2598));
  invx g2500(.A(n2304), .O(n2599));
  invx g2501(.A(n1450), .O(n2600));
  invx g2502(.A(n1444), .O(n2601));
  invx g2503(.A(n1972), .O(n2602));
  invx g2504(.A(n192), .O(n2603));
  invx g2505(.A(n2225), .O(n2604));
  invx g2506(.A(n1469), .O(n2605));
  invx g2507(.A(n1467), .O(n2606));
  invx g2508(.A(n1464), .O(n2607));
  invx g2509(.A(n2007), .O(n2608));
  invx g2510(.A(n1967), .O(n2609));
  invx g2511(.A(n1724), .O(n2610));
  invx g2512(.A(n1446), .O(n2611));
  invx g2513(.A(n1966), .O(n2612));
  invx g2514(.A(n176), .O(n2613));
  invx g2515(.A(n1443), .O(n2614));
  invx g2516(.A(n1543), .O(n2615));
  invx g2517(.A(n1478), .O(n2616));
  invx g2518(.A(n1514), .O(n2617));
  invx g2519(.A(n2087), .O(n2618));
  invx g2520(.A(n1511), .O(n2619));
  invx g2521(.A(n1500), .O(n2620));
  invx g2522(.A(n1501), .O(n2621));
  invx g2523(.A(n1493), .O(n2622));
  invx g2524(.A(n1494), .O(n2623));
  invx g2525(.A(n180), .O(n2624));
  andx g2526(.A(n2626), .B(n2296), .O(n2625));
  andx g2527(.A(n2634), .B(n2627), .O(n2626));
  orx  g2528(.A(n2643), .B(n2628), .O(n2627));
  orx  g2529(.A(n2285), .B(n2629), .O(n2628));
  andx g2530(.A(n2630), .B(n2464), .O(n2629));
  orx  g2531(.A(n2631), .B(n2632), .O(n2630));
  orx  g2532(.A(n2418), .B(n2409), .O(n2631));
  andx g2533(.A(n2319), .B(n2265), .O(n2632));
  invx g2534(.A(pi26), .O(n2633));
  orx  g2535(.A(n2637), .B(n2635), .O(n2634));
  invx g2536(.A(n2636), .O(n2635));
  orx  g2537(.A(n2638), .B(pi32), .O(n2636));
  andx g2538(.A(pi32), .B(n2638), .O(n2637));
  invx g2539(.A(pi33), .O(n2638));
  andx g2540(.A(n1457), .B(n2325), .O(n2639));
  andx g2541(.A(n1455), .B(n2323), .O(n2640));
  andx g2542(.A(n1452), .B(n2310), .O(n2641));
  andx g2543(.A(n2296), .B(n2643), .O(n2642));
  orx  g2544(.A(n2650), .B(n2644), .O(n2643));
  andx g2545(.A(n2645), .B(pi25), .O(n2644));
  andx g2546(.A(n2649), .B(n2646), .O(n2645));
  andx g2547(.A(n2647), .B(pi28), .O(n2646));
  invx g2548(.A(n2648), .O(n2647));
  orx  g2549(.A(n2672), .B(pi26), .O(n2648));
  andx g2550(.A(pi29), .B(pi30), .O(n2649));
  andx g2551(.A(n2652), .B(n2651), .O(n2650));
  invx g2552(.A(pi25), .O(n2651));
  orx  g2553(.A(n2666), .B(n2653), .O(n2652));
  andx g2554(.A(n2654), .B(pi26), .O(n2653));
  orx  g2555(.A(n2655), .B(n2662), .O(n2654));
  andx g2556(.A(n2656), .B(n2402), .O(n2655));
  orx  g2557(.A(n2429), .B(n2657), .O(n2656));
  orx  g2558(.A(n2659), .B(n2658), .O(n2657));
  andx g2559(.A(n2661), .B(n2293), .O(n2658));
  andx g2560(.A(n2660), .B(pi29), .O(n2659));
  invx g2561(.A(n2661), .O(n2660));
  andx g2562(.A(pi31), .B(pi27), .O(n2661));
  andx g2563(.A(n2663), .B(n2292), .O(n2662));
  orx  g2564(.A(n2431), .B(n2664), .O(n2663));
  andx g2565(.A(n2665), .B(pi31), .O(n2664));
  andx g2566(.A(pi30), .B(n2334), .O(n2665));
  andx g2567(.A(n2670), .B(n2667), .O(n2666));
  andx g2568(.A(n2403), .B(n2443), .O(n2667));
  invx g2569(.A(pi28), .O(n2668));
  invx g2570(.A(pi30), .O(n2669));
  andx g2571(.A(n2672), .B(n2671), .O(n2670));
  invx g2572(.A(pi29), .O(n2671));
  andx g2573(.A(n2321), .B(n2353), .O(n2672));
  invx g2574(.A(pi27), .O(n2673));
  andx g2575(.A(n1554), .B(n2311), .O(n2674));
  andx g2576(.A(n1552), .B(n2298), .O(n2675));
  andx g2577(.A(n1550), .B(n2324), .O(n2676));
  andx g2578(.A(n1547), .B(n2309), .O(n2677));
  andx g2579(.A(n1545), .B(n2310), .O(n2678));
  andx g2580(.A(n1540), .B(n2726), .O(n2679));
  andx g2581(.A(n1537), .B(n2325), .O(n2680));
  andx g2582(.A(n1534), .B(n2323), .O(n2681));
  andx g2583(.A(n1531), .B(n2309), .O(n2682));
  andx g2584(.A(n1527), .B(n2311), .O(n2683));
  andx g2585(.A(n1525), .B(n2298), .O(n2684));
  andx g2586(.A(n1523), .B(n2324), .O(n2685));
  andx g2587(.A(n1520), .B(n2323), .O(n2686));
  andx g2588(.A(n1516), .B(n2310), .O(n2687));
  andx g2589(.A(n1513), .B(n2726), .O(n2688));
  andx g2590(.A(n1509), .B(n2325), .O(n2689));
  andx g2591(.A(n1505), .B(n2324), .O(n2690));
  andx g2592(.A(n1498), .B(n2309), .O(n2691));
  andx g2593(.A(n1491), .B(n2311), .O(n2692));
  andx g2594(.A(n1485), .B(n2298), .O(n2693));
  andx g2595(.A(n335), .B(n2325), .O(n2694));
  andx g2596(.A(n333), .B(n2323), .O(n2695));
  andx g2597(.A(n331), .B(n2310), .O(n2696));
  andx g2598(.A(n328), .B(n2296), .O(n2697));
  andx g2599(.A(n325), .B(n2296), .O(n2698));
  andx g2600(.A(n323), .B(n2324), .O(n2699));
  andx g2601(.A(n321), .B(n2309), .O(n2700));
  andx g2602(.A(n315), .B(n2311), .O(n2701));
  andx g2603(.A(n311), .B(n2296), .O(n2702));
  andx g2604(.A(n309), .B(n2325), .O(n2703));
  andx g2605(.A(n305), .B(n2323), .O(n2704));
  andx g2606(.A(n303), .B(n2310), .O(n2705));
  andx g2607(.A(n299), .B(n2311), .O(n2706));
  andx g2608(.A(n295), .B(n2298), .O(n2707));
  andx g2609(.A(n293), .B(n2324), .O(n2708));
  andx g2610(.A(n286), .B(n2309), .O(n2709));
  andx g2611(.A(n282), .B(n2310), .O(n2710));
  andx g2612(.A(n279), .B(n2296), .O(n2711));
  andx g2613(.A(n276), .B(n2325), .O(n2712));
  andx g2614(.A(n272), .B(n2323), .O(n2713));
  andx g2615(.A(n270), .B(n2309), .O(n2714));
  andx g2616(.A(n267), .B(n2311), .O(n2715));
  andx g2617(.A(n263), .B(n2298), .O(n2716));
  andx g2618(.A(n260), .B(n2324), .O(n2717));
  andx g2619(.A(n255), .B(n2323), .O(n2718));
  andx g2620(.A(n249), .B(n2310), .O(n2719));
  andx g2621(.A(n245), .B(n2726), .O(n2720));
  andx g2622(.A(n241), .B(n2325), .O(n2721));
  andx g2623(.A(n232), .B(n2324), .O(n2722));
  andx g2624(.A(n226), .B(n2309), .O(n2723));
  andx g2625(.A(n223), .B(n2311), .O(n2724));
  andx g2626(.A(n217), .B(n2298), .O(n2725));
  invx g2627(.A(n2727), .O(n2726));
  orx  g2628(.A(n2739), .B(n2728), .O(n2727));
  orx  g2629(.A(n2734), .B(n2729), .O(n2728));
  orx  g2630(.A(n2732), .B(n2730), .O(n2729));
  orx  g2631(.A(pi03), .B(n2731), .O(n2730));
  orx  g2632(.A(pi05), .B(pi04), .O(n2731));
  orx  g2633(.A(pi06), .B(n2733), .O(n2732));
  orx  g2634(.A(pi08), .B(pi07), .O(n2733));
  orx  g2635(.A(n2737), .B(n2735), .O(n2734));
  orx  g2636(.A(pi09), .B(n2736), .O(n2735));
  orx  g2637(.A(pi11), .B(pi10), .O(n2736));
  orx  g2638(.A(pi12), .B(n2738), .O(n2737));
  orx  g2639(.A(pi14), .B(pi13), .O(n2738));
  orx  g2640(.A(n2745), .B(n2740), .O(n2739));
  orx  g2641(.A(n2743), .B(n2741), .O(n2740));
  orx  g2642(.A(pi15), .B(n2742), .O(n2741));
  orx  g2643(.A(pi17), .B(pi16), .O(n2742));
  orx  g2644(.A(pi18), .B(n2744), .O(n2743));
  orx  g2645(.A(pi20), .B(pi19), .O(n2744));
  orx  g2646(.A(n2748), .B(n2746), .O(n2745));
  orx  g2647(.A(pi21), .B(n2747), .O(n2746));
  orx  g2648(.A(pi23), .B(pi22), .O(n2747));
  orx  g2649(.A(n2750), .B(n2749), .O(n2748));
  orx  g2650(.A(pi00), .B(pi24), .O(n2749));
  orx  g2651(.A(pi02), .B(pi01), .O(n2750));
endmodule


