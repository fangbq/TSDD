// Benchmark "top" written by ABC on Fri Feb  7 13:27:18 2014

module top ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63;
  wire n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
    n308, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548, n549, n550, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n656, n657,
    n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n669, n670,
    n671, n672, n673, n674, n677, n678, n679, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n729,
    n730, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n745,
    n746, n748, n749, n750, n751, n752, n753, n754, n755, n757, n759, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n813, n814, n817, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n866,
    n867, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1082, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1106, n1107;
  andx g000(.a(pi054), .b(pi056), .O(n297));
  andx g001(.a(n297), .b(pi036), .O(n298));
  invx g002(.a(pi054), .O(n299));
  andx g003(.a(n299), .b(pi056), .O(n300));
  andx g004(.a(n300), .b(pi035), .O(n301));
  orx  g005(.a(n301), .b(n298), .O(n302));
  invx g006(.a(pi056), .O(n303));
  andx g007(.a(n299), .b(n303), .O(n304));
  andx g008(.a(n304), .b(pi037), .O(n305));
  andx g009(.a(pi054), .b(n303), .O(n306));
  andx g010(.a(n306), .b(pi033), .O(n307));
  orx  g011(.a(n307), .b(n305), .O(n308));
  orx  g012(.a(n308), .b(n302), .O(po14));
  andx g013(.a(po14), .b(pi066), .O(n310));
  invx g014(.a(pi066), .O(n311));
  andx g015(.a(n297), .b(pi014), .O(n312));
  andx g016(.a(n300), .b(pi015), .O(n313));
  orx  g017(.a(n313), .b(n312), .O(n314));
  andx g018(.a(n304), .b(pi016), .O(n315));
  andx g019(.a(n306), .b(pi017), .O(n316));
  orx  g020(.a(n316), .b(n315), .O(n317));
  orx  g021(.a(n317), .b(n314), .O(n318));
  andx g022(.a(n318), .b(n311), .O(n319));
  orx  g023(.a(n319), .b(n310), .O(po00));
  invx g024(.a(po14), .O(po01));
  andx g025(.a(n297), .b(pi006), .O(n322));
  andx g026(.a(n300), .b(pi009), .O(n323));
  orx  g027(.a(n323), .b(n322), .O(n324));
  andx g028(.a(n304), .b(pi008), .O(n325));
  andx g029(.a(n306), .b(pi010), .O(n326));
  orx  g030(.a(n326), .b(n325), .O(n327));
  orx  g031(.a(n327), .b(n324), .O(n328));
  andx g032(.a(n328), .b(pi012), .O(n329));
  invx g033(.a(pi012), .O(n330));
  invx g034(.a(n328), .O(n331));
  invx g035(.a(n318), .O(n332));
  invx g036(.a(pi005), .O(n333));
  invx g037(.a(n297), .O(n334));
  orx  g038(.a(n334), .b(n333), .O(n335));
  invx g039(.a(pi002), .O(n336));
  invx g040(.a(n300), .O(n337));
  orx  g041(.a(n337), .b(n336), .O(n338));
  andx g042(.a(n338), .b(n335), .O(n339));
  invx g043(.a(pi003), .O(n340));
  invx g044(.a(n304), .O(n341));
  orx  g045(.a(n341), .b(n340), .O(n342));
  invx g046(.a(pi004), .O(n343));
  invx g047(.a(n306), .O(n344));
  orx  g048(.a(n344), .b(n343), .O(n345));
  andx g049(.a(n345), .b(n342), .O(n346));
  andx g050(.a(n346), .b(n339), .O(n347));
  xorx g051(.a(n347), .b(n332), .O(n348));
  orx  g052(.a(n318), .b(pi013), .O(n349));
  xorx g053(.a(n349), .b(n348), .O(n350));
  xorx g054(.a(n350), .b(n331), .O(n351));
  andx g055(.a(n351), .b(n330), .O(n352));
  orx  g056(.a(n352), .b(n329), .O(po02));
  invx g057(.a(pi049), .O(n354));
  andx g058(.a(n297), .b(pi050), .O(n355));
  andx g059(.a(n300), .b(pi055), .O(n356));
  orx  g060(.a(n356), .b(n355), .O(n357));
  invx g061(.a(n357), .O(n358));
  invx g062(.a(pi052), .O(n359));
  orx  g063(.a(n341), .b(n359), .O(n360));
  andx g064(.a(n306), .b(pi058), .O(n361));
  invx g065(.a(n361), .O(n362));
  andx g066(.a(n362), .b(n360), .O(n363));
  andx g067(.a(n363), .b(n358), .O(po30));
  invx g068(.a(po30), .O(po52));
  andx g069(.a(po52), .b(pi064), .O(n366));
  invx g070(.a(pi064), .O(n367));
  andx g071(.a(pi063), .b(n367), .O(n368));
  orx  g072(.a(n368), .b(n366), .O(n369));
  invx g073(.a(n369), .O(n370));
  andx g074(.a(n370), .b(n354), .O(n371));
  andx g075(.a(n369), .b(pi049), .O(n372));
  invx g076(.a(pi029), .O(n373));
  invx g077(.a(pi028), .O(n374));
  orx  g078(.a(n334), .b(n374), .O(n375));
  invx g079(.a(pi031), .O(n376));
  orx  g080(.a(n337), .b(n376), .O(n377));
  andx g081(.a(n377), .b(n375), .O(n378));
  invx g082(.a(pi030), .O(n379));
  orx  g083(.a(n341), .b(n379), .O(n380));
  invx g084(.a(pi032), .O(n381));
  orx  g085(.a(n344), .b(n381), .O(n382));
  andx g086(.a(n382), .b(n380), .O(n383));
  andx g087(.a(n383), .b(n378), .O(n384));
  orx  g088(.a(n384), .b(n367), .O(n385));
  andx g089(.a(pi000), .b(n367), .O(n386));
  invx g090(.a(n386), .O(n387));
  andx g091(.a(n387), .b(n385), .O(n388));
  andx g092(.a(n388), .b(n373), .O(n389));
  orx  g093(.a(n389), .b(n372), .O(n390));
  orx  g094(.a(n390), .b(n371), .O(n391));
  andx g095(.a(po14), .b(pi064), .O(n392));
  andx g096(.a(pi022), .b(n367), .O(n393));
  orx  g097(.a(n393), .b(n392), .O(n394));
  andx g098(.a(n394), .b(pi034), .O(n395));
  invx g099(.a(n395), .O(n396));
  andx g100(.a(n318), .b(pi064), .O(n397));
  andx g101(.a(pi011), .b(n367), .O(n398));
  orx  g102(.a(n398), .b(n397), .O(n399));
  orx  g103(.a(n399), .b(pi020), .O(n400));
  andx g104(.a(n400), .b(n396), .O(n401));
  orx  g105(.a(n388), .b(n373), .O(n402));
  orx  g106(.a(n394), .b(pi034), .O(n403));
  andx g107(.a(n403), .b(n402), .O(n404));
  andx g108(.a(n404), .b(n401), .O(n405));
  invx g109(.a(n405), .O(n406));
  invx g110(.a(pi019), .O(n407));
  orx  g111(.a(n347), .b(n367), .O(n408));
  andx g112(.a(pi001), .b(n367), .O(n409));
  invx g113(.a(n409), .O(n410));
  andx g114(.a(n410), .b(n408), .O(n411));
  orx  g115(.a(n411), .b(n407), .O(n412));
  invx g116(.a(n412), .O(n413));
  invx g117(.a(pi072), .O(n414));
  andx g118(.a(pi104), .b(pi105), .O(n415));
  andx g119(.a(n415), .b(pi084), .O(n416));
  invx g120(.a(pi104), .O(n417));
  andx g121(.a(n417), .b(pi105), .O(n418));
  andx g122(.a(n418), .b(pi086), .O(n419));
  orx  g123(.a(n419), .b(n416), .O(n420));
  invx g124(.a(n420), .O(n421));
  invx g125(.a(pi077), .O(n422));
  orx  g126(.a(pi104), .b(pi105), .O(n423));
  orx  g127(.a(n423), .b(n422), .O(n424));
  invx g128(.a(pi105), .O(n425));
  andx g129(.a(pi104), .b(n425), .O(n426));
  andx g130(.a(n426), .b(pi080), .O(n427));
  invx g131(.a(n427), .O(n428));
  andx g132(.a(n428), .b(n424), .O(n429));
  andx g133(.a(n429), .b(n421), .O(n430));
  invx g134(.a(n430), .O(n431));
  andx g135(.a(n431), .b(pi123), .O(n432));
  invx g136(.a(pi123), .O(n433));
  andx g137(.a(pi073), .b(n433), .O(n434));
  orx  g138(.a(n434), .b(n432), .O(n435));
  invx g139(.a(n435), .O(n436));
  andx g140(.a(n436), .b(n414), .O(n437));
  orx  g141(.a(n437), .b(n413), .O(n438));
  andx g142(.a(n399), .b(pi020), .O(n439));
  andx g143(.a(n411), .b(n407), .O(n440));
  orx  g144(.a(n440), .b(n439), .O(n441));
  orx  g145(.a(n441), .b(n438), .O(n442));
  orx  g146(.a(n442), .b(n406), .O(n443));
  orx  g147(.a(n443), .b(n391), .O(n444));
  andx g148(.a(n415), .b(pi103), .O(n445));
  andx g149(.a(n418), .b(pi109), .O(n446));
  orx  g150(.a(n446), .b(n445), .O(n447));
  andx g151(.a(n417), .b(n425), .O(n448));
  andx g152(.a(n448), .b(pi101), .O(n449));
  andx g153(.a(n426), .b(pi117), .O(n450));
  orx  g154(.a(n450), .b(n449), .O(n451));
  orx  g155(.a(n451), .b(n447), .O(n452));
  andx g156(.a(n452), .b(pi123), .O(n453));
  andx g157(.a(pi126), .b(n433), .O(n454));
  orx  g158(.a(n454), .b(n453), .O(n455));
  andx g159(.a(n455), .b(pi113), .O(n456));
  invx g160(.a(n456), .O(n457));
  andx g161(.a(n415), .b(pi106), .O(n458));
  andx g162(.a(n418), .b(pi108), .O(n459));
  orx  g163(.a(n459), .b(n458), .O(n460));
  andx g164(.a(n448), .b(pi100), .O(n461));
  andx g165(.a(n426), .b(pi116), .O(n462));
  orx  g166(.a(n462), .b(n461), .O(n463));
  orx  g167(.a(n463), .b(n460), .O(n464));
  andx g168(.a(n464), .b(pi123), .O(n465));
  andx g169(.a(pi124), .b(n433), .O(n466));
  orx  g170(.a(n466), .b(n465), .O(n467));
  andx g171(.a(pi125), .b(pi066), .O(n468));
  andx g172(.a(pi125), .b(n311), .O(n469));
  orx  g173(.a(n469), .b(n468), .O(n470));
  andx g174(.a(n470), .b(n467), .O(n471));
  andx g175(.a(n471), .b(n457), .O(n472));
  andx g176(.a(n415), .b(pi085), .O(n473));
  andx g177(.a(n418), .b(pi089), .O(n474));
  orx  g178(.a(n474), .b(n473), .O(n475));
  invx g179(.a(n475), .O(n476));
  invx g180(.a(pi078), .O(n477));
  orx  g181(.a(n423), .b(n477), .O(n478));
  andx g182(.a(n426), .b(pi081), .O(n479));
  invx g183(.a(n479), .O(n480));
  andx g184(.a(n480), .b(n478), .O(n481));
  andx g185(.a(n481), .b(n476), .O(n482));
  invx g186(.a(n482), .O(n483));
  andx g187(.a(n483), .b(pi123), .O(n484));
  andx g188(.a(pi070), .b(n433), .O(n485));
  orx  g189(.a(n485), .b(n484), .O(n486));
  andx g190(.a(n486), .b(pi067), .O(n487));
  invx g191(.a(n487), .O(n488));
  orx  g192(.a(n455), .b(pi113), .O(n489));
  andx g193(.a(n489), .b(n488), .O(n490));
  andx g194(.a(n415), .b(pi090), .O(n491));
  andx g195(.a(n418), .b(pi087), .O(n492));
  orx  g196(.a(n492), .b(n491), .O(n493));
  invx g197(.a(n493), .O(n494));
  invx g198(.a(pi079), .O(n495));
  orx  g199(.a(n423), .b(n495), .O(n496));
  andx g200(.a(n426), .b(pi082), .O(n497));
  invx g201(.a(n497), .O(n498));
  andx g202(.a(n498), .b(n496), .O(n499));
  andx g203(.a(n499), .b(n494), .O(n500));
  orx  g204(.a(n500), .b(n433), .O(n501));
  andx g205(.a(pi074), .b(n433), .O(n502));
  invx g206(.a(n502), .O(n503));
  andx g207(.a(n503), .b(n501), .O(n504));
  invx g208(.a(n504), .O(n505));
  andx g209(.a(n505), .b(pi083), .O(n506));
  invx g210(.a(n506), .O(n507));
  orx  g211(.a(n486), .b(pi067), .O(n508));
  andx g212(.a(n508), .b(n507), .O(n509));
  andx g213(.a(n509), .b(n490), .O(n510));
  andx g214(.a(n510), .b(n472), .O(n511));
  invx g215(.a(n511), .O(n512));
  andx g216(.a(n415), .b(pi097), .O(n513));
  andx g217(.a(n418), .b(pi095), .O(n514));
  orx  g218(.a(n514), .b(n513), .O(n515));
  andx g219(.a(n448), .b(pi098), .O(n516));
  andx g220(.a(n426), .b(pi096), .O(n517));
  orx  g221(.a(n517), .b(n516), .O(n518));
  orx  g222(.a(n518), .b(n515), .O(n519));
  andx g223(.a(n519), .b(pi123), .O(n520));
  andx g224(.a(pi118), .b(n433), .O(n521));
  orx  g225(.a(n521), .b(n520), .O(n522));
  andx g226(.a(n522), .b(pi094), .O(n523));
  invx g227(.a(n523), .O(n524));
  andx g228(.a(n415), .b(pi091), .O(n525));
  andx g229(.a(n418), .b(pi110), .O(n526));
  orx  g230(.a(n526), .b(n525), .O(n527));
  invx g231(.a(n527), .O(n528));
  invx g232(.a(pi076), .O(n529));
  orx  g233(.a(n423), .b(n529), .O(n530));
  andx g234(.a(n426), .b(pi119), .O(n531));
  invx g235(.a(n531), .O(n532));
  andx g236(.a(n532), .b(n530), .O(n533));
  andx g237(.a(n533), .b(n528), .O(n534));
  invx g238(.a(n534), .O(n535));
  andx g239(.a(n535), .b(pi123), .O(n536));
  andx g240(.a(pi068), .b(n433), .O(n537));
  orx  g241(.a(n537), .b(n536), .O(n538));
  orx  g242(.a(n538), .b(pi038), .O(n539));
  andx g243(.a(n539), .b(n524), .O(n540));
  invx g244(.a(n540), .O(n541));
  andx g245(.a(n297), .b(pi047), .O(n542));
  andx g246(.a(n300), .b(pi044), .O(n543));
  orx  g247(.a(n543), .b(n542), .O(n544));
  invx g248(.a(n544), .O(n545));
  invx g249(.a(pi045), .O(n546));
  orx  g250(.a(n341), .b(n546), .O(n547));
  andx g251(.a(n306), .b(pi048), .O(n548));
  invx g252(.a(n548), .O(n549));
  andx g253(.a(n549), .b(n547), .O(n550));
  andx g254(.a(n550), .b(n545), .O(po59));
  invx g255(.a(po59), .O(po35));
  andx g256(.a(po35), .b(pi064), .O(n553));
  andx g257(.a(pi060), .b(n367), .O(n554));
  orx  g258(.a(n554), .b(n553), .O(n555));
  andx g259(.a(n555), .b(pi046), .O(n556));
  orx  g260(.a(n522), .b(pi094), .O(n557));
  invx g261(.a(n557), .O(n558));
  orx  g262(.a(n558), .b(n556), .O(n559));
  orx  g263(.a(n559), .b(n541), .O(n560));
  andx g264(.a(n415), .b(pi102), .O(n561));
  andx g265(.a(n418), .b(pi092), .O(n562));
  orx  g266(.a(n562), .b(n561), .O(n563));
  andx g267(.a(n448), .b(pi099), .O(n564));
  andx g268(.a(n426), .b(pi093), .O(n565));
  orx  g269(.a(n565), .b(n564), .O(n566));
  orx  g270(.a(n566), .b(n563), .O(n567));
  andx g271(.a(n567), .b(pi123), .O(n568));
  andx g272(.a(pi069), .b(n433), .O(n569));
  orx  g273(.a(n569), .b(n568), .O(n570));
  andx g274(.a(n570), .b(pi039), .O(n571));
  invx g275(.a(pi083), .O(n572));
  andx g276(.a(n504), .b(n572), .O(n573));
  orx  g277(.a(n573), .b(n571), .O(n574));
  andx g278(.a(n538), .b(pi038), .O(n575));
  orx  g279(.a(n570), .b(pi039), .O(n576));
  invx g280(.a(n576), .O(n577));
  orx  g281(.a(n577), .b(n575), .O(n578));
  orx  g282(.a(n578), .b(n574), .O(n579));
  orx  g283(.a(n579), .b(n560), .O(n580));
  andx g284(.a(n297), .b(pi051), .O(n581));
  andx g285(.a(n300), .b(pi057), .O(n582));
  orx  g286(.a(n582), .b(n581), .O(n583));
  andx g287(.a(n304), .b(pi053), .O(n584));
  andx g288(.a(n306), .b(pi059), .O(n585));
  orx  g289(.a(n585), .b(n584), .O(n586));
  orx  g290(.a(n586), .b(n583), .O(po49));
  andx g291(.a(po49), .b(pi064), .O(n588));
  andx g292(.a(pi065), .b(n367), .O(n589));
  orx  g293(.a(n589), .b(n588), .O(n590));
  andx g294(.a(n590), .b(pi062), .O(n591));
  invx g295(.a(n591), .O(n592));
  andx g296(.a(n297), .b(pi025), .O(n593));
  andx g297(.a(n300), .b(pi023), .O(n594));
  orx  g298(.a(n594), .b(n593), .O(n595));
  invx g299(.a(n595), .O(n596));
  invx g300(.a(pi024), .O(n597));
  orx  g301(.a(n341), .b(n597), .O(n598));
  andx g302(.a(n306), .b(pi026), .O(n599));
  invx g303(.a(n599), .O(n600));
  andx g304(.a(n600), .b(n598), .O(n601));
  andx g305(.a(n601), .b(n596), .O(n602));
  invx g306(.a(n602), .O(po50));
  andx g307(.a(po50), .b(pi064), .O(n604));
  andx g308(.a(pi018), .b(n367), .O(n605));
  orx  g309(.a(n605), .b(n604), .O(n606));
  orx  g310(.a(n606), .b(pi027), .O(n607));
  andx g311(.a(n607), .b(n592), .O(n608));
  invx g312(.a(n608), .O(n609));
  andx g313(.a(n435), .b(pi072), .O(n610));
  orx  g314(.a(n590), .b(pi062), .O(n611));
  invx g315(.a(n611), .O(n612));
  orx  g316(.a(n612), .b(n610), .O(n613));
  orx  g317(.a(n613), .b(n609), .O(n614));
  andx g318(.a(n300), .b(pi042), .O(n615));
  orx  g319(.a(n615), .b(n306), .O(n616));
  andx g320(.a(n304), .b(pi040), .O(n617));
  andx g321(.a(n297), .b(pi041), .O(n618));
  orx  g322(.a(n618), .b(n617), .O(n619));
  orx  g323(.a(n619), .b(n616), .O(po13));
  andx g324(.a(po13), .b(pi064), .O(n621));
  andx g325(.a(pi007), .b(n367), .O(n622));
  orx  g326(.a(n622), .b(n621), .O(n623));
  andx g327(.a(n623), .b(pi043), .O(n624));
  invx g328(.a(n624), .O(n625));
  orx  g329(.a(n555), .b(pi046), .O(n626));
  andx g330(.a(n626), .b(n625), .O(n627));
  invx g331(.a(n627), .O(n628));
  andx g332(.a(n606), .b(pi027), .O(n629));
  orx  g333(.a(n623), .b(pi043), .O(n630));
  invx g334(.a(n630), .O(n631));
  orx  g335(.a(n631), .b(n629), .O(n632));
  orx  g336(.a(n632), .b(n628), .O(n633));
  orx  g337(.a(n633), .b(n614), .O(n634));
  orx  g338(.a(n634), .b(n580), .O(n635));
  orx  g339(.a(n635), .b(n512), .O(n636));
  orx  g340(.a(n636), .b(n444), .O(po03));
  andx g341(.a(pi127), .b(pi130), .O(n638));
  andx g342(.a(pi129), .b(pi128), .O(n639));
  andx g343(.a(n639), .b(n638), .O(n640));
  invx g344(.a(n640), .O(n641));
  andx g345(.a(n641), .b(pi131), .O(n642));
  andx g346(.a(pi134), .b(pi133), .O(n643));
  andx g347(.a(pi136), .b(pi135), .O(n644));
  andx g348(.a(n644), .b(n643), .O(n645));
  invx g349(.a(n645), .O(n646));
  andx g350(.a(n646), .b(pi132), .O(n647));
  orx  g351(.a(n647), .b(n642), .O(n648));
  andx g352(.a(pi143), .b(pi144), .O(n649));
  invx g353(.a(pi141), .O(n650));
  invx g354(.a(pi137), .O(n651));
  orx  g355(.a(n651), .b(n650), .O(n652));
  orx  g356(.a(n652), .b(n649), .O(n653));
  orx  g357(.a(n653), .b(n648), .O(po04));
  invx g358(.a(pi135), .O(po05));
  invx g359(.a(n444), .O(n656));
  invx g360(.a(n559), .O(n657));
  andx g361(.a(n657), .b(n540), .O(n658));
  invx g362(.a(n579), .O(n659));
  andx g363(.a(n659), .b(n658), .O(n660));
  invx g364(.a(n613), .O(n661));
  andx g365(.a(n661), .b(n608), .O(n662));
  invx g366(.a(n632), .O(n663));
  andx g367(.a(n663), .b(n627), .O(n664));
  andx g368(.a(n664), .b(n662), .O(n665));
  andx g369(.a(n665), .b(n660), .O(n666));
  andx g370(.a(n666), .b(n511), .O(n667));
  andx g371(.a(n667), .b(n656), .O(po06));
  invx g372(.a(pi038), .O(n669));
  invx g373(.a(pi094), .O(n670));
  orx  g374(.a(n670), .b(n669), .O(n671));
  invx g375(.a(pi039), .O(n672));
  invx g376(.a(pi113), .O(n673));
  orx  g377(.a(n673), .b(n672), .O(n674));
  orx  g378(.a(n674), .b(n671), .O(po07));
  invx g379(.a(pi130), .O(po08));
  invx g380(.a(pi140), .O(n677));
  invx g381(.a(pi139), .O(n678));
  orx  g382(.a(n678), .b(n651), .O(n679));
  orx  g383(.a(n679), .b(n677), .O(po09));
  invx g384(.a(n384), .O(po10));
  invx g385(.a(pi097), .O(n682));
  orx  g386(.a(n417), .b(n425), .O(n683));
  orx  g387(.a(n683), .b(n682), .O(n684));
  invx g388(.a(pi095), .O(n685));
  orx  g389(.a(pi104), .b(n425), .O(n686));
  orx  g390(.a(n686), .b(n685), .O(n687));
  andx g391(.a(n687), .b(n684), .O(n688));
  invx g392(.a(pi098), .O(n689));
  orx  g393(.a(n423), .b(n689), .O(n690));
  invx g394(.a(pi096), .O(n691));
  orx  g395(.a(n417), .b(pi105), .O(n692));
  orx  g396(.a(n692), .b(n691), .O(n693));
  andx g397(.a(n693), .b(n690), .O(n694));
  andx g398(.a(n694), .b(n688), .O(po11));
  invx g399(.a(pi133), .O(po16));
  andx g400(.a(n645), .b(n640), .O(po57));
  invx g401(.a(po57), .O(po17));
  invx g402(.a(pi129), .O(po18));
  invx g403(.a(n648), .O(po19));
  xorx g404(.a(po13), .b(po59), .O(n701));
  xorx g405(.a(n602), .b(po49), .O(n702));
  xorx g406(.a(n702), .b(n701), .O(n703));
  invx g407(.a(n703), .O(n704));
  xorx g408(.a(n384), .b(n318), .O(n705));
  xorx g409(.a(n347), .b(n328), .O(n706));
  xorx g410(.a(po30), .b(po14), .O(n707));
  invx g411(.a(n707), .O(n708));
  andx g412(.a(n708), .b(n706), .O(n709));
  andx g413(.a(n709), .b(n705), .O(n710));
  invx g414(.a(n706), .O(n711));
  andx g415(.a(n707), .b(n705), .O(n712));
  andx g416(.a(n712), .b(n711), .O(n713));
  orx  g417(.a(n713), .b(n710), .O(n714));
  orx  g418(.a(n707), .b(n706), .O(n715));
  orx  g419(.a(n715), .b(n705), .O(n716));
  invx g420(.a(n716), .O(n717));
  invx g421(.a(n705), .O(n718));
  andx g422(.a(n707), .b(n718), .O(n719));
  andx g423(.a(n719), .b(n706), .O(n720));
  orx  g424(.a(n720), .b(n717), .O(n721));
  orx  g425(.a(n721), .b(n714), .O(n722));
  andx g426(.a(n722), .b(n704), .O(n723));
  invx g427(.a(n723), .O(n724));
  invx g428(.a(pi088), .O(n725));
  orx  g429(.a(n722), .b(n704), .O(n726));
  andx g430(.a(n726), .b(n725), .O(n727));
  andx g431(.a(n727), .b(n724), .O(po22));
  andx g432(.a(n318), .b(pi012), .O(n729));
  andx g433(.a(n349), .b(n330), .O(n730));
  orx  g434(.a(n730), .b(n729), .O(po23));
  invx g435(.a(pi134), .O(po24));
  invx g436(.a(pi102), .O(n733));
  orx  g437(.a(n683), .b(n733), .O(n734));
  invx g438(.a(pi092), .O(n735));
  orx  g439(.a(n686), .b(n735), .O(n736));
  andx g440(.a(n736), .b(n734), .O(n737));
  invx g441(.a(pi099), .O(n738));
  orx  g442(.a(n423), .b(n738), .O(n739));
  invx g443(.a(pi093), .O(n740));
  orx  g444(.a(n692), .b(n740), .O(n741));
  andx g445(.a(n741), .b(n739), .O(n742));
  andx g446(.a(n742), .b(n737), .O(po26));
  invx g447(.a(pi114), .O(po28));
  andx g448(.a(po52), .b(pi066), .O(n745));
  andx g449(.a(po10), .b(n311), .O(n746));
  orx  g450(.a(n746), .b(n745), .O(po29));
  andx g451(.a(n464), .b(pi114), .O(n748));
  invx g452(.a(pi114), .O(n749));
  invx g453(.a(n464), .O(n750));
  andx g454(.a(n750), .b(n749), .O(n751));
  andx g455(.a(n692), .b(n423), .O(n752));
  andx g456(.a(n752), .b(n425), .O(n753));
  xorx g457(.a(n753), .b(pi112), .O(n754));
  orx  g458(.a(n754), .b(n751), .O(n755));
  orx  g459(.a(n755), .b(n748), .O(po31));
  invx g460(.a(n347), .O(n757));
  orx  g461(.a(n757), .b(n330), .O(po33));
  invx g462(.a(pi138), .O(n759));
  orx  g463(.a(n759), .b(n651), .O(po34));
  orx  g464(.a(n705), .b(n349), .O(n761));
  orx  g465(.a(n761), .b(n711), .O(n762));
  invx g466(.a(n349), .O(n763));
  orx  g467(.a(n718), .b(n763), .O(n764));
  orx  g468(.a(n764), .b(n711), .O(n765));
  andx g469(.a(n765), .b(n762), .O(n766));
  orx  g470(.a(n705), .b(n763), .O(n767));
  orx  g471(.a(n767), .b(n706), .O(n768));
  orx  g472(.a(n718), .b(n349), .O(n769));
  orx  g473(.a(n769), .b(n706), .O(n770));
  andx g474(.a(n770), .b(n768), .O(n771));
  andx g475(.a(n771), .b(n766), .O(n772));
  xorx g476(.a(n772), .b(n704), .O(n773));
  andx g477(.a(n773), .b(pi066), .O(n774));
  andx g478(.a(n328), .b(n311), .O(n775));
  orx  g479(.a(n775), .b(n774), .O(po36));
  xorx g480(.a(po11), .b(n452), .O(n777));
  xorx g481(.a(n464), .b(n777), .O(n778));
  invx g482(.a(n778), .O(n779));
  xorx g483(.a(n500), .b(n483), .O(n780));
  invx g484(.a(pi107), .O(n781));
  orx  g485(.a(n683), .b(n781), .O(n782));
  invx g486(.a(pi111), .O(n783));
  orx  g487(.a(n686), .b(n783), .O(n784));
  andx g488(.a(n784), .b(n782), .O(n785));
  invx g489(.a(pi075), .O(n786));
  orx  g490(.a(n423), .b(n786), .O(n787));
  invx g491(.a(pi120), .O(n788));
  orx  g492(.a(n692), .b(n788), .O(n789));
  andx g493(.a(n789), .b(n787), .O(n790));
  andx g494(.a(n790), .b(n785), .O(n791));
  xorx g495(.a(n791), .b(n431), .O(n792));
  xorx g496(.a(n567), .b(n534), .O(n793));
  invx g497(.a(n793), .O(n794));
  andx g498(.a(n794), .b(n792), .O(n795));
  andx g499(.a(n795), .b(n780), .O(n796));
  invx g500(.a(n792), .O(n797));
  andx g501(.a(n793), .b(n780), .O(n798));
  andx g502(.a(n798), .b(n797), .O(n799));
  orx  g503(.a(n799), .b(n796), .O(n800));
  orx  g504(.a(n793), .b(n792), .O(n801));
  orx  g505(.a(n801), .b(n780), .O(n802));
  orx  g506(.a(n794), .b(n780), .O(n803));
  orx  g507(.a(n803), .b(n797), .O(n804));
  andx g508(.a(n804), .b(n802), .O(n805));
  invx g509(.a(n805), .O(n806));
  orx  g510(.a(n806), .b(n800), .O(n807));
  andx g511(.a(n807), .b(n779), .O(n808));
  invx g512(.a(n808), .O(n809));
  orx  g513(.a(n807), .b(n779), .O(n810));
  andx g514(.a(n810), .b(n725), .O(n811));
  andx g515(.a(n811), .b(n809), .O(po38));
  andx g516(.a(n349), .b(pi066), .O(n813));
  andx g517(.a(n757), .b(n311), .O(n814));
  orx  g518(.a(n814), .b(n813), .O(po39));
  andx g519(.a(pi146), .b(pi145), .O(po40));
  invx g520(.a(pi132), .O(n817));
  orx  g521(.a(po34), .b(n817), .O(po41));
  xorx g522(.a(pi062), .b(pi027), .O(n819));
  invx g523(.a(pi067), .O(n820));
  xorx g524(.a(pi072), .b(n820), .O(n821));
  xorx g525(.a(n821), .b(n819), .O(n822));
  invx g526(.a(pi034), .O(n823));
  xorx g527(.a(pi049), .b(n823), .O(n824));
  invx g528(.a(n824), .O(n825));
  xorx g529(.a(pi071), .b(n373), .O(n826));
  invx g530(.a(n826), .O(n827));
  invx g531(.a(pi043), .O(n828));
  xorx g532(.a(pi046), .b(n828), .O(n829));
  orx  g533(.a(n829), .b(n827), .O(n830));
  orx  g534(.a(n830), .b(n825), .O(n831));
  invx g535(.a(n829), .O(n832));
  orx  g536(.a(n832), .b(n825), .O(n833));
  orx  g537(.a(n833), .b(n826), .O(n834));
  andx g538(.a(n834), .b(n831), .O(n835));
  orx  g539(.a(n829), .b(n826), .O(n836));
  orx  g540(.a(n836), .b(n824), .O(n837));
  orx  g541(.a(n832), .b(n824), .O(n838));
  orx  g542(.a(n838), .b(n827), .O(n839));
  andx g543(.a(n839), .b(n837), .O(n840));
  andx g544(.a(n840), .b(n835), .O(n841));
  xorx g545(.a(n841), .b(n822), .O(n842));
  invx g546(.a(n842), .O(po42));
  invx g547(.a(n452), .O(po45));
  xorx g548(.a(pi112), .b(n749), .O(n845));
  xorx g549(.a(pi038), .b(n672), .O(n846));
  invx g550(.a(n846), .O(n847));
  xorx g551(.a(pi115), .b(n572), .O(n848));
  invx g552(.a(n848), .O(n849));
  xorx g553(.a(pi113), .b(n670), .O(n850));
  orx  g554(.a(n850), .b(n849), .O(n851));
  orx  g555(.a(n851), .b(n847), .O(n852));
  invx g556(.a(n850), .O(n853));
  orx  g557(.a(n853), .b(n847), .O(n854));
  orx  g558(.a(n854), .b(n848), .O(n855));
  andx g559(.a(n855), .b(n852), .O(n856));
  orx  g560(.a(n850), .b(n848), .O(n857));
  orx  g561(.a(n857), .b(n846), .O(n858));
  orx  g562(.a(n853), .b(n846), .O(n859));
  orx  g563(.a(n859), .b(n849), .O(n860));
  andx g564(.a(n860), .b(n858), .O(n861));
  andx g565(.a(n861), .b(n856), .O(n862));
  xorx g566(.a(n862), .b(n845), .O(n863));
  invx g567(.a(n863), .O(po46));
  invx g568(.a(pi127), .O(po47));
  invx g569(.a(pi142), .O(n866));
  orx  g570(.a(n652), .b(n866), .O(n867));
  orx  g571(.a(n867), .b(n648), .O(po48));
  invx g572(.a(pi122), .O(n869));
  andx g573(.a(n567), .b(n869), .O(n870));
  andx g574(.a(po11), .b(pi121), .O(n871));
  andx g575(.a(n871), .b(n870), .O(n872));
  orx  g576(.a(n872), .b(pi020), .O(n873));
  orx  g577(.a(po26), .b(pi122), .O(n874));
  invx g578(.a(pi121), .O(n875));
  orx  g579(.a(n519), .b(n875), .O(n876));
  orx  g580(.a(n876), .b(n874), .O(n877));
  orx  g581(.a(n877), .b(pi083), .O(n878));
  andx g582(.a(n878), .b(n873), .O(n879));
  xorx g583(.a(n879), .b(n332), .O(n880));
  invx g584(.a(n880), .O(n881));
  orx  g585(.a(n872), .b(pi029), .O(n882));
  orx  g586(.a(n877), .b(pi038), .O(n883));
  andx g587(.a(n883), .b(n882), .O(n884));
  xorx g588(.a(n884), .b(po10), .O(n885));
  andx g589(.a(n877), .b(n407), .O(n886));
  andx g590(.a(n872), .b(n820), .O(n887));
  orx  g591(.a(n887), .b(n886), .O(n888));
  andx g592(.a(n888), .b(n347), .O(n889));
  andx g593(.a(n889), .b(n885), .O(n890));
  andx g594(.a(n890), .b(n881), .O(n891));
  orx  g595(.a(n884), .b(po10), .O(n892));
  invx g596(.a(n892), .O(n893));
  invx g597(.a(pi020), .O(n894));
  andx g598(.a(n877), .b(n894), .O(n895));
  andx g599(.a(n872), .b(n572), .O(n896));
  orx  g600(.a(n896), .b(n895), .O(n897));
  andx g601(.a(n897), .b(n332), .O(n898));
  andx g602(.a(n898), .b(n885), .O(n899));
  orx  g603(.a(n899), .b(n893), .O(n900));
  orx  g604(.a(n900), .b(n891), .O(n901));
  andx g605(.a(po35), .b(pi061), .O(n902));
  invx g606(.a(n902), .O(n903));
  invx g607(.a(pi046), .O(n904));
  andx g608(.a(n877), .b(n904), .O(n905));
  andx g609(.a(n872), .b(n673), .O(n906));
  orx  g610(.a(n906), .b(n905), .O(n907));
  andx g611(.a(n907), .b(pi061), .O(n908));
  xorx g612(.a(n908), .b(n903), .O(n909));
  andx g613(.a(po52), .b(pi061), .O(n910));
  invx g614(.a(n910), .O(n911));
  andx g615(.a(n877), .b(n354), .O(n912));
  andx g616(.a(n872), .b(n670), .O(n913));
  orx  g617(.a(n913), .b(n912), .O(n914));
  andx g618(.a(n914), .b(pi061), .O(n915));
  xorx g619(.a(n915), .b(n911), .O(n916));
  orx  g620(.a(n872), .b(pi034), .O(n917));
  orx  g621(.a(n877), .b(pi039), .O(n918));
  andx g622(.a(n918), .b(n917), .O(n919));
  xorx g623(.a(n919), .b(po14), .O(n920));
  andx g624(.a(po13), .b(pi061), .O(n921));
  invx g625(.a(n921), .O(n922));
  orx  g626(.a(n922), .b(n872), .O(n923));
  andx g627(.a(pi061), .b(n828), .O(n924));
  andx g628(.a(n924), .b(n877), .O(n925));
  xorx g629(.a(n925), .b(n923), .O(n926));
  andx g630(.a(po49), .b(pi061), .O(n927));
  invx g631(.a(n927), .O(n928));
  orx  g632(.a(n928), .b(n872), .O(n929));
  invx g633(.a(pi062), .O(n930));
  andx g634(.a(pi061), .b(n930), .O(n931));
  andx g635(.a(n931), .b(n877), .O(n932));
  xorx g636(.a(n932), .b(n929), .O(n933));
  andx g637(.a(n933), .b(n926), .O(n934));
  andx g638(.a(n934), .b(n920), .O(n935));
  andx g639(.a(n935), .b(n916), .O(n936));
  andx g640(.a(n936), .b(n909), .O(n937));
  andx g641(.a(n937), .b(n901), .O(n938));
  andx g642(.a(n877), .b(n823), .O(n939));
  andx g643(.a(n872), .b(n672), .O(n940));
  orx  g644(.a(n940), .b(n939), .O(n941));
  andx g645(.a(n941), .b(po01), .O(n942));
  andx g646(.a(n942), .b(n926), .O(n943));
  andx g647(.a(n943), .b(n933), .O(n944));
  andx g648(.a(n944), .b(n909), .O(n945));
  andx g649(.a(n945), .b(n916), .O(n946));
  andx g650(.a(n915), .b(n911), .O(n947));
  andx g651(.a(n947), .b(n934), .O(n948));
  andx g652(.a(n948), .b(n909), .O(n949));
  andx g653(.a(n908), .b(n903), .O(n950));
  andx g654(.a(n950), .b(n934), .O(n951));
  andx g655(.a(n932), .b(n929), .O(n952));
  andx g656(.a(n925), .b(n923), .O(n953));
  andx g657(.a(n953), .b(n933), .O(n954));
  orx  g658(.a(n954), .b(n952), .O(n955));
  orx  g659(.a(n955), .b(n951), .O(n956));
  orx  g660(.a(n956), .b(n949), .O(n957));
  orx  g661(.a(n957), .b(n946), .O(n958));
  orx  g662(.a(n958), .b(n938), .O(n959));
  andx g663(.a(n871), .b(n874), .O(n960));
  invx g664(.a(n960), .O(n961));
  orx  g665(.a(n872), .b(n500), .O(n962));
  orx  g666(.a(n962), .b(n961), .O(n963));
  andx g667(.a(n877), .b(n572), .O(n964));
  andx g668(.a(n964), .b(n960), .O(n965));
  xorx g669(.a(n965), .b(n963), .O(n966));
  orx  g670(.a(n872), .b(n602), .O(n967));
  orx  g671(.a(n967), .b(n961), .O(n968));
  invx g672(.a(pi027), .O(n969));
  andx g673(.a(n877), .b(n969), .O(n970));
  andx g674(.a(n970), .b(n960), .O(n971));
  xorx g675(.a(n971), .b(n968), .O(n972));
  andx g676(.a(n972), .b(n966), .O(n973));
  orx  g677(.a(n872), .b(n482), .O(n974));
  orx  g678(.a(n974), .b(n961), .O(n975));
  andx g679(.a(n877), .b(n820), .O(n976));
  andx g680(.a(n976), .b(n960), .O(n977));
  xorx g681(.a(n977), .b(n975), .O(n978));
  orx  g682(.a(n872), .b(n430), .O(n979));
  orx  g683(.a(n979), .b(n961), .O(n980));
  andx g684(.a(n877), .b(n414), .O(n981));
  andx g685(.a(n981), .b(n960), .O(n982));
  xorx g686(.a(n982), .b(n980), .O(n983));
  andx g687(.a(n983), .b(n978), .O(n984));
  andx g688(.a(n984), .b(n973), .O(n985));
  andx g689(.a(n982), .b(n980), .O(n986));
  andx g690(.a(n986), .b(n966), .O(n987));
  andx g691(.a(n987), .b(n978), .O(n988));
  andx g692(.a(n971), .b(n968), .O(n989));
  andx g693(.a(n989), .b(n978), .O(n990));
  andx g694(.a(n983), .b(n966), .O(n991));
  andx g695(.a(n991), .b(n990), .O(n992));
  andx g696(.a(n965), .b(n963), .O(n993));
  andx g697(.a(n977), .b(n975), .O(n994));
  andx g698(.a(n994), .b(n966), .O(n995));
  orx  g699(.a(n995), .b(n993), .O(n996));
  orx  g700(.a(n996), .b(n992), .O(n997));
  orx  g701(.a(n997), .b(n988), .O(n998));
  orx  g702(.a(n998), .b(n985), .O(n999));
  andx g703(.a(n999), .b(n959), .O(n1000));
  xorx g704(.a(n884), .b(n384), .O(n1001));
  orx  g705(.a(n872), .b(pi019), .O(n1002));
  orx  g706(.a(n877), .b(pi067), .O(n1003));
  andx g707(.a(n1003), .b(n1002), .O(n1004));
  orx  g708(.a(n1004), .b(n757), .O(n1005));
  orx  g709(.a(n1005), .b(n1001), .O(n1006));
  orx  g710(.a(n1006), .b(n880), .O(n1007));
  orx  g711(.a(n879), .b(n318), .O(n1008));
  orx  g712(.a(n1008), .b(n1001), .O(n1009));
  andx g713(.a(n1009), .b(n892), .O(n1010));
  andx g714(.a(n1010), .b(n1007), .O(n1011));
  xorx g715(.a(n908), .b(n902), .O(n1012));
  xorx g716(.a(n915), .b(n910), .O(n1013));
  xorx g717(.a(n919), .b(po01), .O(n1014));
  andx g718(.a(n921), .b(n877), .O(n1015));
  xorx g719(.a(n925), .b(n1015), .O(n1016));
  andx g720(.a(n927), .b(n877), .O(n1017));
  xorx g721(.a(n932), .b(n1017), .O(n1018));
  orx  g722(.a(n1018), .b(n1016), .O(n1019));
  orx  g723(.a(n1019), .b(n1014), .O(n1020));
  orx  g724(.a(n1020), .b(n1013), .O(n1021));
  orx  g725(.a(n1021), .b(n1012), .O(n1022));
  orx  g726(.a(n1022), .b(n1011), .O(n1023));
  orx  g727(.a(n919), .b(po14), .O(n1024));
  orx  g728(.a(n1024), .b(n1016), .O(n1025));
  orx  g729(.a(n1025), .b(n1018), .O(n1026));
  orx  g730(.a(n1026), .b(n1012), .O(n1027));
  orx  g731(.a(n1027), .b(n1013), .O(n1028));
  invx g732(.a(pi061), .O(n1029));
  orx  g733(.a(n872), .b(pi049), .O(n1030));
  orx  g734(.a(n877), .b(pi094), .O(n1031));
  andx g735(.a(n1031), .b(n1030), .O(n1032));
  orx  g736(.a(n1032), .b(n1029), .O(n1033));
  orx  g737(.a(n1033), .b(n910), .O(n1034));
  orx  g738(.a(n1034), .b(n1019), .O(n1035));
  orx  g739(.a(n1035), .b(n1012), .O(n1036));
  orx  g740(.a(n872), .b(pi046), .O(n1037));
  orx  g741(.a(n877), .b(pi113), .O(n1038));
  andx g742(.a(n1038), .b(n1037), .O(n1039));
  orx  g743(.a(n1039), .b(n1029), .O(n1040));
  orx  g744(.a(n1040), .b(n902), .O(n1041));
  orx  g745(.a(n1041), .b(n1019), .O(n1042));
  invx g746(.a(n952), .O(n1043));
  invx g747(.a(n924), .O(n1044));
  orx  g748(.a(n1044), .b(n872), .O(n1045));
  orx  g749(.a(n1045), .b(n1015), .O(n1046));
  orx  g750(.a(n1046), .b(n1018), .O(n1047));
  andx g751(.a(n1047), .b(n1043), .O(n1048));
  andx g752(.a(n1048), .b(n1042), .O(n1049));
  andx g753(.a(n1049), .b(n1036), .O(n1050));
  andx g754(.a(n1050), .b(n1028), .O(n1051));
  andx g755(.a(n1051), .b(n1023), .O(n1052));
  andx g756(.a(n998), .b(n1052), .O(n1053));
  orx  g757(.a(n1053), .b(n1000), .O(po51));
  xorx g758(.a(pi150), .b(pi149), .O(n1055));
  xorx g759(.a(pi019), .b(n894), .O(n1056));
  xorx g760(.a(n1056), .b(n1055), .O(n1057));
  xorx g761(.a(pi156), .b(pi155), .O(n1058));
  invx g762(.a(n1058), .O(n1059));
  xorx g763(.a(pi152), .b(pi151), .O(n1060));
  invx g764(.a(n1060), .O(n1061));
  xorx g765(.a(pi154), .b(pi153), .O(n1062));
  andx g766(.a(n1062), .b(n1061), .O(n1063));
  andx g767(.a(n1063), .b(n1059), .O(n1064));
  invx g768(.a(n1062), .O(n1065));
  andx g769(.a(n1065), .b(n1059), .O(n1066));
  andx g770(.a(n1066), .b(n1060), .O(n1067));
  orx  g771(.a(n1067), .b(n1064), .O(n1068));
  andx g772(.a(n1062), .b(n1060), .O(n1069));
  andx g773(.a(n1069), .b(n1058), .O(n1070));
  andx g774(.a(n1065), .b(n1058), .O(n1071));
  andx g775(.a(n1071), .b(n1061), .O(n1072));
  orx  g776(.a(n1072), .b(n1070), .O(n1073));
  orx  g777(.a(n1073), .b(n1068), .O(n1074));
  andx g778(.a(n1074), .b(n1057), .O(n1075));
  invx g779(.a(n1075), .O(n1076));
  orx  g780(.a(n1074), .b(n1057), .O(n1077));
  andx g781(.a(n1077), .b(pi021), .O(n1078));
  andx g782(.a(n1078), .b(n1076), .O(po54));
  invx g783(.a(pi128), .O(po55));
  invx g784(.a(pi136), .O(po58));
  invx g785(.a(pi131), .O(n1082));
  orx  g786(.a(po34), .b(n1082), .O(po61));
  invx g787(.a(n800), .O(n1084));
  andx g788(.a(n805), .b(n1084), .O(n1085));
  andx g789(.a(n1085), .b(n778), .O(n1086));
  orx  g790(.a(n1086), .b(pi088), .O(n1087));
  orx  g791(.a(n1087), .b(n808), .O(n1088));
  orx  g792(.a(n707), .b(n711), .O(n1089));
  orx  g793(.a(n1089), .b(n718), .O(n1090));
  invx g794(.a(n713), .O(n1091));
  andx g795(.a(n1091), .b(n1090), .O(n1092));
  orx  g796(.a(n708), .b(n705), .O(n1093));
  orx  g797(.a(n1093), .b(n711), .O(n1094));
  andx g798(.a(n1094), .b(n716), .O(n1095));
  andx g799(.a(n1095), .b(n1092), .O(n1096));
  andx g800(.a(n1096), .b(n703), .O(n1097));
  orx  g801(.a(n1097), .b(pi088), .O(n1098));
  orx  g802(.a(n1098), .b(n723), .O(n1099));
  invx g803(.a(po54), .O(n1100));
  andx g804(.a(n842), .b(po19), .O(n1101));
  andx g805(.a(n1101), .b(n863), .O(n1102));
  andx g806(.a(n1102), .b(n1100), .O(n1103));
  andx g807(.a(n1103), .b(n1099), .O(n1104));
  andx g808(.a(n1104), .b(n1088), .O(po62));
  invx g809(.a(n1103), .O(n1106));
  orx  g810(.a(n1106), .b(po22), .O(n1107));
  orx  g811(.a(n1107), .b(po38), .O(po63));
  bufx g812(.a(pi148), .O(po12));
  bufx g813(.a(pi147), .O(po15));
  orx  g814(.a(n319), .b(n310), .O(po20));
  bufx g815(.a(pi145), .O(po21));
  bufx g816(.a(pi148), .O(po25));
  bufx g817(.a(pi147), .O(po27));
  bufx g818(.a(pi147), .O(po32));
  bufx g819(.a(pi145), .O(po37));
  orx  g820(.a(n746), .b(n745), .O(po43));
  bufx g821(.a(pi145), .O(po44));
  orx  g822(.a(n775), .b(n774), .O(po53));
  orx  g823(.a(n814), .b(n813), .O(po56));
  bufx g824(.a(pi145), .O(po60));
endmodule


